module __sobel_filter__sobel_filter_4(
  input wire [511:0] in_img,
  (*keep*) output wire [127:0] out
);
  // lint_off MULTIPLY
  function automatic [47:0] umul48b_24b_x_24b (input reg [23:0] lhs, input reg [23:0] rhs);
    begin
      umul48b_24b_x_24b = lhs * rhs;
    end
  endfunction
  // lint_on MULTIPLY
  wire [31:0] in_img_unflattened[16];
  assign in_img_unflattened[0] = in_img[31:0];
  assign in_img_unflattened[1] = in_img[63:32];
  assign in_img_unflattened[2] = in_img[95:64];
  assign in_img_unflattened[3] = in_img[127:96];
  assign in_img_unflattened[4] = in_img[159:128];
  assign in_img_unflattened[5] = in_img[191:160];
  assign in_img_unflattened[6] = in_img[223:192];
  assign in_img_unflattened[7] = in_img[255:224];
  assign in_img_unflattened[8] = in_img[287:256];
  assign in_img_unflattened[9] = in_img[319:288];
  assign in_img_unflattened[10] = in_img[351:320];
  assign in_img_unflattened[11] = in_img[383:352];
  assign in_img_unflattened[12] = in_img[415:384];
  assign in_img_unflattened[13] = in_img[447:416];
  assign in_img_unflattened[14] = in_img[479:448];
  assign in_img_unflattened[15] = in_img[511:480];
  wire [31:0] array_index_157912;
  wire [31:0] array_index_157913;
  wire [31:0] array_index_157914;
  wire [31:0] array_index_157915;
  wire result_sign__389;
  wire [7:0] x_bexp__73;
  wire result_sign__482;
  wire [7:0] x_bexp__145;
  wire result_sign__579;
  wire [7:0] x_bexp__289;
  wire result_sign__681;
  wire [7:0] x_bexp__433;
  wire result_sign__390;
  wire [8:0] add_157933;
  wire [7:0] x_bexp__664;
  wire result_sign__94;
  wire [22:0] x_fraction__73;
  wire result_sign__483;
  wire [8:0] add_157938;
  wire [7:0] x_bexp__665;
  wire result_sign__481;
  wire [22:0] x_fraction__145;
  wire result_sign__580;
  wire [8:0] add_157943;
  wire [7:0] x_bexp__666;
  wire result_sign__578;
  wire [22:0] x_fraction__289;
  wire result_sign__682;
  wire [8:0] add_157948;
  wire [7:0] x_bexp__667;
  wire result_sign__680;
  wire [22:0] x_fraction__433;
  wire ne_157954;
  wire ne_157959;
  wire ne_157964;
  wire ne_157969;
  wire [9:0] exp__36;
  wire [23:0] x_fraction__74;
  wire [9:0] exp__83;
  wire [9:0] sign_ext_157977;
  wire [23:0] x_fraction__147;
  wire [9:0] exp__165;
  wire [9:0] sign_ext_157981;
  wire [23:0] x_fraction__291;
  wire [9:0] exp__246;
  wire [9:0] sign_ext_157985;
  wire [23:0] x_fraction__435;
  wire [9:0] exp__37;
  wire [23:0] x_fraction__75;
  wire result_sign__796;
  wire result_sign__797;
  wire [9:0] exp__85;
  wire [23:0] x_fraction__149;
  wire result_sign__798;
  wire result_sign__799;
  wire [9:0] exp__167;
  wire [23:0] x_fraction__293;
  wire result_sign__800;
  wire result_sign__801;
  wire [9:0] exp__248;
  wire [23:0] x_fraction__437;
  wire result_sign__802;
  wire result_sign__803;
  wire [24:0] concat_158012;
  wire [24:0] concat_158013;
  wire [24:0] concat_158015;
  wire [24:0] concat_158016;
  wire [24:0] concat_158018;
  wire [24:0] concat_158019;
  wire [24:0] sel_158020;
  wire [24:0] sel_158021;
  wire [24:0] sel_158022;
  wire [24:0] sel_158023;
  wire result_sign__928;
  wire [22:0] fraction__86;
  wire result_sign__934;
  wire [22:0] fraction__190;
  wire result_sign__940;
  wire [22:0] fraction__369;
  wire result_sign__948;
  wire [22:0] fraction__548;
  wire [23:0] fraction__87;
  wire [23:0] fraction__192;
  wire [23:0] fraction__371;
  wire [23:0] fraction__550;
  wire do_round_up__18;
  wire [23:0] add_158049;
  wire do_round_up__40;
  wire [23:0] add_158051;
  wire do_round_up__79;
  wire [23:0] add_158053;
  wire do_round_up__118;
  wire [23:0] add_158055;
  wire [23:0] fraction__88;
  wire [23:0] fraction__194;
  wire [23:0] fraction__373;
  wire [23:0] fraction__552;
  wire [9:0] add_158065;
  wire [9:0] add_158067;
  wire [9:0] add_158069;
  wire [9:0] add_158071;
  wire [9:0] exp__39;
  wire [9:0] exp__89;
  wire [9:0] exp__171;
  wire [9:0] exp__253;
  wire [8:0] result_exp__27;
  wire [8:0] result_exp__61;
  wire [8:0] result_exp__121;
  wire [8:0] result_exp__181;
  wire [7:0] high_exp__9;
  wire [22:0] result_fraction__8;
  wire [8:0] result_exp__28;
  wire [7:0] high_exp__143;
  wire [22:0] result_fraction__543;
  wire [8:0] result_exp__63;
  wire [7:0] high_exp__209;
  wire [22:0] result_fraction__610;
  wire [8:0] result_exp__123;
  wire [7:0] high_exp__277;
  wire [22:0] result_fraction__677;
  wire [8:0] result_exp__183;
  wire eq_158104;
  wire is_result_nan__3;
  wire is_result_nan__24;
  wire is_result_nan__84;
  wire has_inf_arg__9;
  wire and_reduce_158122;
  wire is_subnormal__9;
  wire [22:0] result_fraction__481;
  wire has_inf_arg__21;
  wire and_reduce_158127;
  wire is_subnormal__21;
  wire [22:0] result_fraction__544;
  wire has_inf_arg__41;
  wire and_reduce_158132;
  wire is_subnormal__41;
  wire [22:0] result_fraction__611;
  wire has_inf_arg__61;
  wire and_reduce_158137;
  wire is_subnormal__61;
  wire [22:0] result_fraction__678;
  wire ne_158141;
  wire ne_158143;
  wire ne_158145;
  wire ne_158147;
  wire is_result_nan__18;
  wire is_result_nan__40;
  wire is_result_nan__79;
  wire is_result_nan__118;
  wire [22:0] result_fraction__54;
  wire or_158158;
  wire [7:0] high_exp__81;
  wire [22:0] result_fraction__118;
  wire or_158162;
  wire [7:0] high_exp__144;
  wire [22:0] result_fraction__235;
  wire or_158166;
  wire [7:0] high_exp__210;
  wire [22:0] result_fraction__352;
  wire or_158170;
  wire [7:0] high_exp__278;
  wire [22:0] result_fraction__55;
  wire [22:0] nan_fraction__9;
  wire [7:0] result_exp__29;
  wire [7:0] x_bexp__668;
  wire [22:0] result_fraction__120;
  wire [22:0] nan_fraction__107;
  wire [7:0] result_exp__65;
  wire [7:0] x_bexp__669;
  wire [22:0] result_fraction__237;
  wire [22:0] nan_fraction__134;
  wire [7:0] result_exp__125;
  wire [7:0] x_bexp__670;
  wire [22:0] result_fraction__354;
  wire [22:0] nan_fraction__163;
  wire [7:0] result_exp__185;
  wire [7:0] x_bexp__671;
  wire [22:0] result_fraction__56;
  wire [22:0] result_fraction__122;
  wire [22:0] result_fraction__239;
  wire [22:0] result_fraction__356;
  wire [27:0] wide_x__18;
  wire [27:0] wide_x__39;
  wire [27:0] wide_x__77;
  wire [27:0] wide_x__115;
  wire x_sign__19;
  wire [27:0] wide_x__19;
  wire x_sign__37;
  wire [27:0] wide_x__41;
  wire x_sign__73;
  wire [27:0] wide_x__79;
  wire x_sign__109;
  wire [27:0] wide_x__117;
  wire result_sign__45;
  wire [27:0] neg_158222;
  wire result_sign__98;
  wire [27:0] neg_158225;
  wire result_sign__195;
  wire [27:0] neg_158228;
  wire result_sign__292;
  wire [27:0] neg_158231;
  wire result_sign__46;
  wire result_sign__100;
  wire result_sign__197;
  wire result_sign__294;
  wire [24:0] sel_158244;
  wire [24:0] sel_158246;
  wire [24:0] sel_158248;
  wire [24:0] sel_158250;
  wire [27:0] xddend_x__10;
  wire [27:0] xddend_x__19;
  wire [27:0] xddend_x__37;
  wire [27:0] xddend_x__55;
  wire [28:0] fraction__89;
  wire [27:0] neg_158257;
  wire [28:0] fraction__196;
  wire [27:0] neg_158259;
  wire [28:0] fraction__375;
  wire [27:0] neg_158261;
  wire [28:0] fraction__554;
  wire [27:0] neg_158263;
  wire result_sign__47;
  wire result_sign__102;
  wire result_sign__199;
  wire result_sign__296;
  wire [24:0] sel_158272;
  wire [24:0] sel_158273;
  wire [24:0] sel_158274;
  wire [24:0] sel_158275;
  wire [27:0] concat_158284;
  wire [27:0] concat_158285;
  wire [27:0] concat_158286;
  wire [27:0] concat_158287;
  wire [28:0] one_hot_158288;
  wire [28:0] one_hot_158289;
  wire [28:0] one_hot_158290;
  wire [28:0] one_hot_158291;
  wire [4:0] encode_158292;
  wire [4:0] encode_158293;
  wire [4:0] encode_158294;
  wire [4:0] encode_158295;
  wire [22:0] result_fraction__482;
  wire [22:0] result_fraction__545;
  wire [22:0] result_fraction__612;
  wire [22:0] result_fraction__679;
  wire cancel__10;
  wire carry_bit__9;
  wire [27:0] leading_zeroes__9;
  wire cancel__20;
  wire carry_bit__20;
  wire [27:0] leading_zeroes__20;
  wire [31:0] array_index_158318;
  wire cancel__39;
  wire carry_bit__39;
  wire [27:0] leading_zeroes__39;
  wire cancel__58;
  wire carry_bit__58;
  wire [27:0] leading_zeroes__58;
  wire [31:0] array_index_158331;
  wire [27:0] add_158335;
  wire [27:0] add_158339;
  wire [7:0] x_bexp__157;
  wire [27:0] add_158344;
  wire [27:0] add_158348;
  wire [7:0] x_bexp__445;
  wire [26:0] cancel_fraction__9;
  wire result_sign__956;
  wire [26:0] cancel_fraction__20;
  wire result_sign__957;
  wire [26:0] cancel_fraction__39;
  wire result_sign__958;
  wire [26:0] cancel_fraction__58;
  wire result_sign__959;
  wire [2:0] concat_158374;
  wire [2:0] concat_158379;
  wire [2:0] concat_158384;
  wire [2:0] concat_158389;
  wire result_sign__960;
  wire [23:0] one_hot_sel_158396;
  wire result_sign__1104;
  wire [1:0] add_158398;
  wire result_sign__961;
  wire [23:0] one_hot_sel_158402;
  wire result_sign__1106;
  wire [1:0] add_158404;
  wire [7:0] x_bexp__672;
  wire result_sign__484;
  wire [22:0] x_fraction__157;
  wire result_sign__962;
  wire [23:0] one_hot_sel_158411;
  wire result_sign__1108;
  wire [1:0] add_158413;
  wire result_sign__963;
  wire [23:0] one_hot_sel_158417;
  wire result_sign__1112;
  wire [1:0] add_158419;
  wire [7:0] x_bexp__673;
  wire result_sign__683;
  wire [22:0] x_fraction__445;
  wire ne_158434;
  wire ne_158447;
  wire nor_158451;
  wire result_sign__1116;
  wire [24:0] add_158453;
  wire [9:0] exp__40;
  wire nor_158456;
  wire result_sign__1117;
  wire [24:0] add_158458;
  wire [9:0] exp__91;
  wire [9:0] sign_ext_158460;
  wire [23:0] x_fraction__159;
  wire nor_158464;
  wire result_sign__1118;
  wire [24:0] add_158466;
  wire [9:0] exp__173;
  wire nor_158469;
  wire result_sign__1119;
  wire [24:0] add_158471;
  wire [9:0] exp__255;
  wire [9:0] sign_ext_158473;
  wire [23:0] x_fraction__447;
  wire do_round_up__19;
  wire [9:0] exp__41;
  wire do_round_up__42;
  wire [9:0] exp__93;
  wire [23:0] x_fraction__161;
  wire result_sign__804;
  wire result_sign__805;
  wire do_round_up__81;
  wire [9:0] exp__175;
  wire do_round_up__120;
  wire [9:0] exp__257;
  wire [23:0] x_fraction__449;
  wire result_sign__806;
  wire result_sign__807;
  wire [25:0] sel_158502;
  wire [25:0] sel_158504;
  wire [24:0] concat_158506;
  wire [24:0] concat_158507;
  wire [25:0] sel_158508;
  wire [25:0] sel_158510;
  wire [24:0] concat_158512;
  wire [24:0] concat_158513;
  wire result_sign__391;
  wire [7:0] x_bexp__648;
  wire rounding_carry__9;
  wire [24:0] sel_158517;
  wire result_sign__486;
  wire [7:0] x_bexp__649;
  wire rounding_carry__20;
  wire [24:0] sel_158521;
  wire result_sign__581;
  wire [7:0] x_bexp__650;
  wire rounding_carry__39;
  wire [24:0] sel_158525;
  wire result_sign__685;
  wire [7:0] x_bexp__651;
  wire rounding_carry__58;
  wire [24:0] sel_158529;
  wire result_sign__929;
  wire [22:0] fraction__95;
  wire result_sign__935;
  wire [22:0] fraction__208;
  wire result_sign__941;
  wire [22:0] fraction__387;
  wire result_sign__949;
  wire [22:0] fraction__566;
  wire result_sign__392;
  wire [8:0] add_158547;
  wire [23:0] fraction__96;
  wire result_sign__487;
  wire [8:0] add_158553;
  wire [23:0] fraction__210;
  wire result_sign__582;
  wire [8:0] add_158559;
  wire [23:0] fraction__389;
  wire result_sign__686;
  wire [8:0] add_158565;
  wire [23:0] fraction__568;
  wire do_round_up__20;
  wire [23:0] add_158576;
  wire do_round_up__44;
  wire [23:0] add_158583;
  wire do_round_up__83;
  wire [23:0] add_158590;
  wire do_round_up__122;
  wire [23:0] add_158597;
  wire [9:0] add_158598;
  wire [23:0] fraction__97;
  wire [9:0] add_158603;
  wire [23:0] fraction__212;
  wire [9:0] add_158608;
  wire [23:0] fraction__391;
  wire [9:0] add_158613;
  wire [23:0] fraction__570;
  wire [9:0] wide_exponent__27;
  wire [9:0] add_158621;
  wire [9:0] wide_exponent__58;
  wire [9:0] add_158625;
  wire [9:0] wide_exponent__115;
  wire [9:0] add_158629;
  wire [9:0] wide_exponent__172;
  wire [9:0] add_158633;
  wire [9:0] wide_exponent__28;
  wire [9:0] exp__43;
  wire [9:0] wide_exponent__60;
  wire [9:0] exp__97;
  wire [9:0] wide_exponent__117;
  wire [9:0] exp__179;
  wire [9:0] wide_exponent__174;
  wire [9:0] exp__261;
  wire [8:0] result_exp__30;
  wire [8:0] result_exp__67;
  wire [8:0] result_exp__127;
  wire [8:0] result_exp__187;
  wire [8:0] result_exp__31;
  wire [7:0] high_exp__146;
  wire [22:0] result_fraction__548;
  wire [22:0] result_fraction__547;
  wire [8:0] result_exp__69;
  wire [8:0] result_exp__129;
  wire [7:0] high_exp__280;
  wire [22:0] result_fraction__682;
  wire [22:0] result_fraction__681;
  wire [8:0] result_exp__189;
  wire [8:0] wide_exponent__29;
  wire [22:0] result_fraction__770;
  wire [22:0] result_fraction__483;
  wire [8:0] wide_exponent__62;
  wire [22:0] result_fraction__803;
  wire [22:0] result_fraction__546;
  wire is_result_nan__45;
  wire ne_158692;
  wire [8:0] wide_exponent__119;
  wire [22:0] result_fraction__836;
  wire [22:0] result_fraction__613;
  wire [8:0] wide_exponent__176;
  wire [22:0] result_fraction__869;
  wire [22:0] result_fraction__680;
  wire is_result_nan__123;
  wire ne_158703;
  wire ne_158707;
  wire and_reduce_158711;
  wire ne_158713;
  wire is_result_nan__44;
  wire has_inf_arg__24;
  wire and_reduce_158719;
  wire ne_158721;
  wire and_reduce_158725;
  wire ne_158727;
  wire is_result_nan__122;
  wire has_inf_arg__64;
  wire and_reduce_158733;
  wire is_result_nan__19;
  wire is_operand_inf__9;
  wire and_reduce_158740;
  wire [7:0] high_exp__83;
  wire is_result_nan__42;
  wire is_operand_inf__20;
  wire and_reduce_158749;
  wire [7:0] high_exp__147;
  wire is_result_nan__81;
  wire is_operand_inf__39;
  wire and_reduce_158758;
  wire [7:0] high_exp__212;
  wire is_result_nan__120;
  wire is_operand_inf__58;
  wire and_reduce_158767;
  wire [7:0] high_exp__281;
  wire [2:0] fraction_shift__29;
  wire [2:0] fraction_shift__28;
  wire is_subnormal__10;
  wire [7:0] high_exp__82;
  wire [7:0] result_exp__32;
  wire [2:0] fraction_shift__385;
  wire [2:0] fraction_shift__263;
  wire is_subnormal__23;
  wire [7:0] high_exp__145;
  wire [7:0] result_exp__71;
  wire [2:0] fraction_shift__403;
  wire [2:0] fraction_shift__298;
  wire is_subnormal__43;
  wire [7:0] high_exp__211;
  wire [7:0] result_exp__131;
  wire [2:0] fraction_shift__421;
  wire [2:0] fraction_shift__333;
  wire is_subnormal__63;
  wire [7:0] high_exp__279;
  wire [7:0] result_exp__191;
  wire [7:0] result_exp__6;
  wire [27:0] rounded_fraction__9;
  wire [2:0] fraction_shift__30;
  wire result_sign__393;
  wire [7:0] result_exponent__10;
  wire result_sign__394;
  wire [7:0] result_exp__72;
  wire [27:0] rounded_fraction__20;
  wire [2:0] fraction_shift__62;
  wire result_sign__488;
  wire [7:0] result_exponent__20;
  wire result_sign__489;
  wire [7:0] result_exp__132;
  wire [27:0] rounded_fraction__39;
  wire [2:0] fraction_shift__119;
  wire result_sign__583;
  wire [7:0] result_exponent__39;
  wire result_sign__584;
  wire [7:0] result_exp__192;
  wire [27:0] rounded_fraction__58;
  wire [2:0] fraction_shift__176;
  wire result_sign__687;
  wire [7:0] result_exponent__58;
  wire result_sign__688;
  wire result_sign__395;
  wire [27:0] shrl_158840;
  wire [8:0] concat_158843;
  wire result_sign__490;
  wire [27:0] shrl_158847;
  wire [8:0] concat_158850;
  wire result_sign__585;
  wire [27:0] shrl_158854;
  wire [8:0] concat_158857;
  wire [8:0] concat_158858;
  wire result_sign__689;
  wire [27:0] shrl_158861;
  wire [8:0] concat_158864;
  wire [8:0] concat_158865;
  wire [22:0] result_fraction__57;
  wire [22:0] result_fraction__60;
  wire [8:0] sum__10;
  wire [22:0] result_fraction__124;
  wire [22:0] result_fraction__130;
  wire [8:0] sum__22;
  wire [8:0] concat_158878;
  wire [22:0] result_fraction__241;
  wire [22:0] result_fraction__247;
  wire [8:0] sum__41;
  wire [8:0] concat_158884;
  wire [22:0] result_fraction__358;
  wire [22:0] result_fraction__364;
  wire [8:0] sum__60;
  wire [8:0] sum__2;
  wire [22:0] result_fraction__58;
  wire [22:0] nan_fraction__81;
  wire [22:0] result_fraction__61;
  wire [22:0] nan_fraction__82;
  wire [8:0] sum__23;
  wire [22:0] result_fraction__126;
  wire [22:0] nan_fraction__108;
  wire [22:0] result_fraction__132;
  wire [22:0] nan_fraction__109;
  wire [8:0] sum__42;
  wire [22:0] result_fraction__243;
  wire [22:0] nan_fraction__135;
  wire [22:0] result_fraction__249;
  wire [22:0] nan_fraction__136;
  wire [8:0] sum__61;
  wire [22:0] result_fraction__360;
  wire [22:0] nan_fraction__164;
  wire [22:0] result_fraction__366;
  wire [22:0] nan_fraction__165;
  wire [22:0] result_fraction__59;
  wire [22:0] result_fraction__62;
  wire [7:0] prod_bexp__42;
  wire [7:0] x_bexp__674;
  wire [22:0] result_fraction__128;
  wire [22:0] result_fraction__134;
  wire [7:0] prod_bexp__83;
  wire [7:0] x_bexp__675;
  wire [22:0] result_fraction__245;
  wire [22:0] result_fraction__251;
  wire [7:0] prod_bexp__155;
  wire [7:0] x_bexp__676;
  wire [22:0] result_fraction__362;
  wire [22:0] result_fraction__368;
  wire [7:0] prod_bexp__227;
  wire [7:0] x_bexp__677;
  wire [22:0] result_fraction__469;
  wire [7:0] prod_bexp__6;
  wire [7:0] x_bexp__678;
  wire [22:0] prod_fraction__30;
  wire [7:0] incremented_sum__78;
  wire [22:0] result_fraction__470;
  wire [7:0] prod_bexp__84;
  wire [7:0] x_bexp__679;
  wire [22:0] prod_fraction__61;
  wire [7:0] incremented_sum__96;
  wire [22:0] result_fraction__471;
  wire [7:0] prod_bexp__156;
  wire [7:0] x_bexp__680;
  wire [22:0] prod_fraction__115;
  wire [7:0] incremented_sum__114;
  wire [22:0] result_fraction__472;
  wire [7:0] prod_bexp__228;
  wire [7:0] x_bexp__681;
  wire [22:0] prod_fraction__169;
  wire [7:0] incremented_sum__132;
  wire [22:0] prod_fraction__4;
  wire [7:0] incremented_sum__79;
  wire [27:0] wide_y__20;
  wire [7:0] x_bexpbs_difference__11;
  wire [22:0] prod_fraction__62;
  wire [7:0] incremented_sum__97;
  wire [27:0] wide_y__43;
  wire [7:0] x_bexpbs_difference__21;
  wire [22:0] prod_fraction__116;
  wire [7:0] incremented_sum__115;
  wire [27:0] wide_y__81;
  wire [7:0] x_bexpbs_difference__39;
  wire [22:0] prod_fraction__170;
  wire [7:0] incremented_sum__133;
  wire [27:0] wide_y__119;
  wire [7:0] x_bexpbs_difference__57;
  wire [27:0] wide_y__3;
  wire [7:0] x_bexpbs_difference__2;
  wire has_pos_inf__9;
  wire [7:0] x_bexp__86;
  wire [7:0] x_bexp__682;
  wire [27:0] wide_y__21;
  wire [7:0] sub_159038;
  wire [27:0] wide_y__44;
  wire [7:0] x_bexpbs_difference__22;
  wire has_pos_inf__20;
  wire [7:0] x_bexp__171;
  wire [7:0] x_bexp__683;
  wire [27:0] wide_y__45;
  wire [7:0] sub_159047;
  wire [27:0] wide_y__82;
  wire [7:0] x_bexpbs_difference__40;
  wire has_pos_inf__39;
  wire [7:0] x_bexp__315;
  wire [7:0] x_bexp__684;
  wire [27:0] wide_y__83;
  wire [7:0] sub_159056;
  wire [27:0] wide_y__120;
  wire [7:0] x_bexpbs_difference__58;
  wire has_pos_inf__58;
  wire [7:0] x_bexp__459;
  wire [7:0] x_bexp__685;
  wire [27:0] wide_y__121;
  wire [7:0] sub_159065;
  wire [7:0] x_bexp__14;
  wire [7:0] x_bexp__686;
  wire [27:0] wide_y__4;
  wire [7:0] sub_159069;
  wire [22:0] x_fraction__86;
  wire [27:0] dropped__10;
  wire [7:0] x_bexp__172;
  wire [7:0] x_bexp__687;
  wire [27:0] wide_y__46;
  wire [7:0] sub_159079;
  wire x_sign__41;
  wire [22:0] x_fraction__171;
  wire [27:0] dropped__22;
  wire [7:0] x_bexp__316;
  wire [7:0] x_bexp__688;
  wire [27:0] wide_y__84;
  wire [7:0] sub_159090;
  wire [22:0] x_fraction__315;
  wire [27:0] dropped__41;
  wire [7:0] x_bexp__460;
  wire [7:0] x_bexp__689;
  wire [27:0] wide_y__122;
  wire [7:0] sub_159100;
  wire x_sign__113;
  wire [22:0] x_fraction__459;
  wire [27:0] dropped__60;
  wire [7:0] high_exp__479;
  wire [22:0] x_fraction__14;
  wire [27:0] dropped__2;
  wire result_sign__48;
  wire [27:0] wide_x__20;
  wire [7:0] high_exp__481;
  wire [22:0] x_fraction__172;
  wire [27:0] dropped__23;
  wire nand_159126;
  wire result_sign__108;
  wire result_sign__104;
  wire [27:0] wide_x__43;
  wire [7:0] high_exp__483;
  wire [22:0] x_fraction__316;
  wire [27:0] dropped__42;
  wire result_sign__201;
  wire [27:0] wide_x__81;
  wire [7:0] high_exp__486;
  wire [22:0] x_fraction__460;
  wire [27:0] dropped__61;
  wire nand_159152;
  wire result_sign__302;
  wire result_sign__298;
  wire [27:0] wide_x__119;
  wire [27:0] wide_x__3;
  wire result_sign__49;
  wire [27:0] wide_x__21;
  wire [27:0] wide_x__44;
  wire result_sign__110;
  wire result_sign__106;
  wire [27:0] wide_x__45;
  wire [27:0] wide_x__82;
  wire result_sign__203;
  wire [27:0] wide_x__83;
  wire [27:0] wide_x__120;
  wire result_sign__304;
  wire result_sign__300;
  wire [27:0] wide_x__121;
  wire result_sign__7;
  wire [27:0] wide_x__4;
  wire x_sign__22;
  wire prod_sign__10;
  wire [27:0] neg_159204;
  wire [27:0] sticky__32;
  wire result_sign__111;
  wire [27:0] wide_x__46;
  wire x_sign__43;
  wire prod_sign__21;
  wire [27:0] neg_159213;
  wire [27:0] sticky__70;
  wire result_sign__208;
  wire [27:0] wide_x__84;
  wire x_sign__79;
  wire prod_sign__39;
  wire [27:0] neg_159222;
  wire [27:0] sticky__129;
  wire result_sign__305;
  wire [27:0] wide_x__122;
  wire x_sign__115;
  wire prod_sign__57;
  wire [27:0] neg_159231;
  wire [27:0] sticky__188;
  wire x_sign__4;
  wire prod_sign__2;
  wire [27:0] neg_159236;
  wire [27:0] sticky__6;
  wire [27:0] xddend_y__10;
  wire x_sign__44;
  wire prod_sign__22;
  wire [27:0] neg_159245;
  wire [27:0] sticky__71;
  wire [27:0] xddend_y__21;
  wire x_sign__80;
  wire prod_sign__40;
  wire [27:0] neg_159254;
  wire [27:0] sticky__130;
  wire [27:0] xddend_y__39;
  wire x_sign__116;
  wire prod_sign__58;
  wire [27:0] neg_159263;
  wire [27:0] sticky__189;
  wire [27:0] xddend_y__57;
  wire [27:0] xddend_y__2;
  wire [24:0] sel_159274;
  wire result_sign__964;
  wire [27:0] xddend_y__22;
  wire [24:0] sel_159281;
  wire result_sign__965;
  wire [27:0] xddend_y__40;
  wire [24:0] sel_159288;
  wire result_sign__966;
  wire [27:0] xddend_y__58;
  wire [24:0] sel_159295;
  wire result_sign__967;
  wire [24:0] sel_159298;
  wire result_sign__968;
  wire [24:0] sel_159303;
  wire result_sign__969;
  wire [24:0] sel_159308;
  wire result_sign__970;
  wire [24:0] sel_159313;
  wire result_sign__971;
  wire [25:0] add_159320;
  wire [25:0] add_159323;
  wire [25:0] add_159326;
  wire [25:0] add_159329;
  wire [25:0] add_159330;
  wire [25:0] add_159333;
  wire [25:0] add_159336;
  wire [25:0] add_159339;
  wire [27:0] concat_159344;
  wire [27:0] concat_159347;
  wire [27:0] concat_159350;
  wire [27:0] concat_159353;
  wire [27:0] concat_159354;
  wire [27:0] concat_159357;
  wire [27:0] concat_159360;
  wire [27:0] concat_159363;
  wire [27:0] xbs_fraction__10;
  wire [27:0] xbs_fraction__21;
  wire [27:0] xbs_fraction__39;
  wire [27:0] xbs_fraction__57;
  wire [27:0] xbs_fraction__2;
  wire [27:0] reverse_159379;
  wire [27:0] xbs_fraction__22;
  wire [27:0] reverse_159381;
  wire [27:0] xbs_fraction__40;
  wire [27:0] reverse_159383;
  wire [27:0] xbs_fraction__58;
  wire [27:0] reverse_159385;
  wire [27:0] reverse_159386;
  wire [28:0] one_hot_159387;
  wire [27:0] reverse_159388;
  wire [28:0] one_hot_159389;
  wire [27:0] reverse_159390;
  wire [28:0] one_hot_159391;
  wire [27:0] reverse_159392;
  wire [28:0] one_hot_159393;
  wire [28:0] one_hot_159394;
  wire [4:0] encode_159395;
  wire [28:0] one_hot_159396;
  wire [4:0] encode_159397;
  wire [28:0] one_hot_159398;
  wire [4:0] encode_159399;
  wire [28:0] one_hot_159400;
  wire [4:0] encode_159401;
  wire [4:0] encode_159402;
  wire [4:0] encode_159404;
  wire [4:0] encode_159406;
  wire [4:0] encode_159408;
  wire cancel__11;
  wire carry_bit__10;
  wire [22:0] result_fraction__484;
  wire cancel__22;
  wire carry_bit__22;
  wire [22:0] result_fraction__549;
  wire cancel__41;
  wire carry_bit__41;
  wire [22:0] result_fraction__614;
  wire cancel__60;
  wire carry_bit__60;
  wire [22:0] result_fraction__683;
  wire cancel__1;
  wire carry_bit__2;
  wire [22:0] result_fraction__485;
  wire [27:0] leading_zeroes__10;
  wire cancel__23;
  wire carry_bit__23;
  wire [22:0] result_fraction__550;
  wire [27:0] leading_zeroes__22;
  wire cancel__42;
  wire carry_bit__42;
  wire [22:0] result_fraction__615;
  wire [27:0] leading_zeroes__41;
  wire cancel__61;
  wire carry_bit__61;
  wire [22:0] result_fraction__684;
  wire [27:0] leading_zeroes__60;
  wire [27:0] leading_zeroes__2;
  wire [26:0] carry_fraction__20;
  wire [27:0] add_159476;
  wire [27:0] leading_zeroes__23;
  wire [26:0] carry_fraction__43;
  wire [27:0] add_159489;
  wire [31:0] array_index_159490;
  wire [27:0] leading_zeroes__42;
  wire [26:0] carry_fraction__81;
  wire [27:0] add_159503;
  wire [27:0] leading_zeroes__61;
  wire [26:0] carry_fraction__119;
  wire [27:0] add_159516;
  wire [31:0] array_index_159517;
  wire [26:0] carry_fraction__3;
  wire [27:0] add_159524;
  wire [2:0] concat_159525;
  wire [26:0] carry_fraction__21;
  wire [26:0] cancel_fraction__10;
  wire result_sign__485;
  wire [26:0] carry_fraction__44;
  wire [27:0] add_159535;
  wire [2:0] concat_159536;
  wire [26:0] carry_fraction__45;
  wire [26:0] cancel_fraction__22;
  wire result_sign__492;
  wire [7:0] x_bexp__173;
  wire [26:0] carry_fraction__82;
  wire [27:0] add_159547;
  wire [2:0] concat_159548;
  wire [26:0] carry_fraction__83;
  wire [26:0] cancel_fraction__41;
  wire result_sign__684;
  wire [26:0] carry_fraction__120;
  wire [27:0] add_159558;
  wire [2:0] concat_159559;
  wire [26:0] carry_fraction__121;
  wire [26:0] cancel_fraction__60;
  wire result_sign__691;
  wire [7:0] x_bexp__461;
  wire [2:0] concat_159564;
  wire [26:0] carry_fraction__4;
  wire [26:0] cancel_fraction__2;
  wire [26:0] shifted_fraction__10;
  wire [2:0] concat_159570;
  wire [26:0] carry_fraction__46;
  wire [26:0] cancel_fraction__23;
  wire [26:0] shifted_fraction__22;
  wire [2:0] concat_159576;
  wire [26:0] carry_fraction__84;
  wire [26:0] cancel_fraction__42;
  wire [26:0] shifted_fraction__41;
  wire [2:0] concat_159582;
  wire [26:0] carry_fraction__122;
  wire [26:0] cancel_fraction__61;
  wire [26:0] shifted_fraction__60;
  wire [26:0] shifted_fraction__2;
  wire result_sign__972;
  wire result_sign__398;
  wire [8:0] add_159592;
  wire [26:0] shifted_fraction__23;
  wire result_sign__973;
  wire result_sign__495;
  wire [8:0] add_159597;
  wire [7:0] x_bexp__690;
  wire result_sign__491;
  wire [22:0] x_fraction__173;
  wire [26:0] shifted_fraction__42;
  wire result_sign__974;
  wire result_sign__588;
  wire [8:0] add_159605;
  wire [26:0] shifted_fraction__61;
  wire result_sign__975;
  wire result_sign__694;
  wire [8:0] add_159610;
  wire [7:0] x_bexp__691;
  wire result_sign__690;
  wire [22:0] x_fraction__461;
  wire result_sign__976;
  wire [2:0] normal_chunk__10;
  wire [2:0] fraction_shift__229;
  wire [1:0] half_way_chunk__10;
  wire result_sign__977;
  wire [2:0] normal_chunk__22;
  wire [2:0] fraction_shift__264;
  wire [1:0] half_way_chunk__22;
  wire ne_159634;
  wire result_sign__978;
  wire [2:0] normal_chunk__41;
  wire [2:0] fraction_shift__299;
  wire [1:0] half_way_chunk__41;
  wire result_sign__979;
  wire [2:0] normal_chunk__60;
  wire [2:0] fraction_shift__334;
  wire [1:0] half_way_chunk__60;
  wire ne_159657;
  wire [2:0] normal_chunk__2;
  wire [2:0] fraction_shift__230;
  wire [1:0] half_way_chunk__2;
  wire result_sign__396;
  wire [24:0] add_159669;
  wire [9:0] exp__44;
  wire [2:0] normal_chunk__23;
  wire [2:0] fraction_shift__265;
  wire [1:0] half_way_chunk__23;
  wire result_sign__493;
  wire [24:0] add_159680;
  wire [9:0] exp__99;
  wire [23:0] x_fraction__175;
  wire [2:0] normal_chunk__42;
  wire [2:0] fraction_shift__300;
  wire [1:0] half_way_chunk__42;
  wire result_sign__586;
  wire [24:0] add_159694;
  wire [9:0] exp__181;
  wire [2:0] normal_chunk__61;
  wire [2:0] fraction_shift__335;
  wire [1:0] half_way_chunk__61;
  wire result_sign__692;
  wire [24:0] add_159705;
  wire [9:0] exp__263;
  wire [9:0] sign_ext_159707;
  wire [23:0] x_fraction__463;
  wire result_sign__397;
  wire [24:0] add_159713;
  wire do_round_up__21;
  wire [9:0] exp__45;
  wire result_sign__494;
  wire [24:0] add_159722;
  wire do_round_up__46;
  wire [9:0] exp__101;
  wire [23:0] x_fraction__177;
  wire result_sign__808;
  wire result_sign__809;
  wire result_sign__587;
  wire [24:0] add_159734;
  wire do_round_up__85;
  wire [9:0] exp__183;
  wire result_sign__693;
  wire [24:0] add_159743;
  wire do_round_up__124;
  wire [9:0] exp__265;
  wire [23:0] x_fraction__465;
  wire result_sign__810;
  wire result_sign__811;
  wire do_round_up__4;
  wire [27:0] rounded_fraction__10;
  wire do_round_up__47;
  wire [27:0] rounded_fraction__22;
  wire do_round_up__86;
  wire [27:0] rounded_fraction__41;
  wire do_round_up__125;
  wire [27:0] rounded_fraction__60;
  wire [24:0] concat_159774;
  wire [24:0] concat_159775;
  wire [27:0] rounded_fraction__2;
  wire result_sign__399;
  wire [7:0] x_bexp__77;
  wire rounding_carry__10;
  wire [24:0] sel_159780;
  wire [27:0] rounded_fraction__23;
  wire result_sign__496;
  wire [7:0] x_bexp__594;
  wire rounding_carry__22;
  wire [24:0] sel_159785;
  wire [27:0] rounded_fraction__42;
  wire result_sign__589;
  wire [7:0] x_bexp__612;
  wire rounding_carry__41;
  wire [24:0] sel_159790;
  wire [27:0] rounded_fraction__61;
  wire result_sign__695;
  wire [7:0] x_bexp__630;
  wire rounding_carry__60;
  wire [24:0] sel_159795;
  wire result_sign__400;
  wire [7:0] x_bexp__577;
  wire rounding_carry__2;
  wire result_sign__930;
  wire [22:0] fraction__104;
  wire result_sign__497;
  wire [7:0] x_bexp__595;
  wire rounding_carry__23;
  wire result_sign__936;
  wire [22:0] fraction__226;
  wire result_sign__590;
  wire [7:0] x_bexp__613;
  wire rounding_carry__42;
  wire result_sign__942;
  wire [22:0] fraction__405;
  wire result_sign__696;
  wire [7:0] x_bexp__631;
  wire rounding_carry__61;
  wire result_sign__950;
  wire [22:0] fraction__584;
  wire result_sign__401;
  wire [8:0] add_159827;
  wire [23:0] fraction__105;
  wire result_sign__498;
  wire [8:0] add_159837;
  wire [23:0] fraction__228;
  wire result_sign__591;
  wire [8:0] add_159847;
  wire [23:0] fraction__407;
  wire result_sign__697;
  wire [8:0] add_159857;
  wire [23:0] fraction__586;
  wire result_sign__402;
  wire [8:0] add_159865;
  wire do_round_up__22;
  wire [23:0] add_159874;
  wire result_sign__499;
  wire [8:0] add_159876;
  wire do_round_up__48;
  wire [23:0] add_159885;
  wire result_sign__592;
  wire [8:0] add_159887;
  wire do_round_up__87;
  wire [23:0] add_159896;
  wire result_sign__698;
  wire [8:0] add_159898;
  wire do_round_up__126;
  wire [23:0] add_159907;
  wire [9:0] add_159913;
  wire [23:0] fraction__106;
  wire [9:0] add_159923;
  wire [23:0] fraction__230;
  wire [9:0] add_159933;
  wire [23:0] fraction__409;
  wire [9:0] add_159943;
  wire [23:0] fraction__588;
  wire [9:0] add_159948;
  wire [9:0] wide_exponent__30;
  wire [9:0] add_159954;
  wire [9:0] add_159955;
  wire [9:0] wide_exponent__64;
  wire [9:0] add_159961;
  wire [9:0] add_159962;
  wire [9:0] wide_exponent__121;
  wire [9:0] add_159968;
  wire [9:0] add_159969;
  wire [9:0] wide_exponent__178;
  wire [9:0] add_159975;
  wire [9:0] wide_exponent__4;
  wire [9:0] wide_exponent__31;
  wire [9:0] exp__47;
  wire [9:0] wide_exponent__65;
  wire [9:0] wide_exponent__66;
  wire [9:0] exp__105;
  wire [9:0] wide_exponent__122;
  wire [9:0] wide_exponent__123;
  wire [9:0] exp__187;
  wire [9:0] wide_exponent__179;
  wire [9:0] wide_exponent__180;
  wire [9:0] exp__269;
  wire [9:0] wide_exponent__5;
  wire [7:0] high_exp__365;
  wire [22:0] result_fraction__771;
  wire [7:0] high_exp__366;
  wire [22:0] result_fraction__772;
  wire [7:0] high_exp__84;
  wire [22:0] result_fraction__486;
  wire [7:0] high_exp__85;
  wire [22:0] result_fraction__487;
  wire [9:0] wide_exponent__67;
  wire [7:0] high_exp__397;
  wire [22:0] result_fraction__804;
  wire [7:0] high_exp__398;
  wire [22:0] result_fraction__805;
  wire [7:0] high_exp__148;
  wire [22:0] result_fraction__551;
  wire [7:0] high_exp__149;
  wire [22:0] result_fraction__552;
  wire [9:0] wide_exponent__124;
  wire [7:0] high_exp__429;
  wire [22:0] result_fraction__837;
  wire [7:0] high_exp__430;
  wire [22:0] result_fraction__838;
  wire [7:0] high_exp__213;
  wire [22:0] result_fraction__616;
  wire [7:0] high_exp__214;
  wire [22:0] result_fraction__617;
  wire [9:0] wide_exponent__181;
  wire [7:0] high_exp__461;
  wire [22:0] result_fraction__870;
  wire [7:0] high_exp__462;
  wire [22:0] result_fraction__871;
  wire [7:0] high_exp__282;
  wire [22:0] result_fraction__685;
  wire [7:0] high_exp__283;
  wire [22:0] result_fraction__686;
  wire ne_160043;
  wire ne_160045;
  wire eq_160046;
  wire eq_160047;
  wire eq_160048;
  wire eq_160049;
  wire [8:0] result_exp__33;
  wire ne_160055;
  wire ne_160057;
  wire eq_160058;
  wire eq_160059;
  wire eq_160060;
  wire eq_160061;
  wire [8:0] result_exp__73;
  wire ne_160067;
  wire ne_160069;
  wire eq_160070;
  wire eq_160071;
  wire eq_160072;
  wire eq_160073;
  wire [8:0] result_exp__133;
  wire ne_160079;
  wire ne_160081;
  wire eq_160082;
  wire eq_160083;
  wire eq_160084;
  wire eq_160085;
  wire [8:0] result_exp__193;
  wire [8:0] result_exp__34;
  wire [7:0] high_exp__153;
  wire [22:0] result_fraction__556;
  wire [22:0] result_fraction__555;
  wire [8:0] result_exp__75;
  wire [8:0] result_exp__135;
  wire [7:0] high_exp__287;
  wire [22:0] result_fraction__690;
  wire [22:0] result_fraction__689;
  wire [8:0] result_exp__195;
  wire [7:0] high_exp__86;
  wire [22:0] result_fraction__756;
  wire [7:0] high_exp__87;
  wire [22:0] result_fraction__757;
  wire [22:0] result_fraction__488;
  wire [22:0] result_fraction__489;
  wire [8:0] wide_exponent__32;
  wire has_pos_inf__10;
  wire has_neg_inf__10;
  wire [7:0] high_exp__150;
  wire [22:0] result_fraction__789;
  wire [7:0] high_exp__151;
  wire [22:0] result_fraction__790;
  wire [22:0] result_fraction__553;
  wire [22:0] result_fraction__554;
  wire [8:0] wide_exponent__68;
  wire has_pos_inf__22;
  wire has_neg_inf__22;
  wire eq_160149;
  wire ne_160150;
  wire [7:0] high_exp__215;
  wire [22:0] result_fraction__822;
  wire [7:0] high_exp__216;
  wire [22:0] result_fraction__823;
  wire [22:0] result_fraction__618;
  wire [22:0] result_fraction__619;
  wire [8:0] wide_exponent__125;
  wire has_pos_inf__41;
  wire has_neg_inf__41;
  wire [7:0] high_exp__284;
  wire [22:0] result_fraction__855;
  wire [7:0] high_exp__285;
  wire [22:0] result_fraction__856;
  wire [22:0] result_fraction__687;
  wire [22:0] result_fraction__688;
  wire [8:0] wide_exponent__182;
  wire has_pos_inf__60;
  wire has_neg_inf__60;
  wire is_result_nan__60;
  wire ne_160177;
  wire [8:0] wide_exponent__6;
  wire eq_160181;
  wire ne_160182;
  wire eq_160183;
  wire ne_160184;
  wire and_reduce_160195;
  wire [8:0] wide_exponent__69;
  wire eq_160197;
  wire ne_160198;
  wire eq_160199;
  wire ne_160200;
  wire is_result_nan__48;
  wire has_inf_arg__25;
  wire and_reduce_160213;
  wire [8:0] wide_exponent__126;
  wire eq_160215;
  wire ne_160216;
  wire eq_160217;
  wire ne_160218;
  wire and_reduce_160229;
  wire [8:0] wide_exponent__183;
  wire eq_160231;
  wire ne_160232;
  wire eq_160233;
  wire ne_160234;
  wire is_result_nan__126;
  wire has_inf_arg__65;
  wire and_reduce_160247;
  wire is_result_nan__21;
  wire is_operand_inf__10;
  wire and_reduce_160260;
  wire [7:0] high_exp__90;
  wire is_result_nan__46;
  wire is_operand_inf__22;
  wire and_reduce_160275;
  wire [7:0] high_exp__155;
  wire is_result_nan__85;
  wire is_operand_inf__41;
  wire and_reduce_160290;
  wire [7:0] high_exp__219;
  wire is_result_nan__124;
  wire is_operand_inf__60;
  wire and_reduce_160305;
  wire [7:0] high_exp__289;
  wire is_result_nan__4;
  wire is_operand_inf__2;
  wire and_reduce_160313;
  wire [2:0] fraction_shift__368;
  wire [2:0] fraction_shift__231;
  wire is_subnormal__11;
  wire [7:0] high_exp__88;
  wire [7:0] result_exp__35;
  wire is_result_nan__47;
  wire is_operand_inf__23;
  wire and_reduce_160326;
  wire [2:0] fraction_shift__386;
  wire [2:0] fraction_shift__266;
  wire is_subnormal__25;
  wire [7:0] high_exp__152;
  wire [7:0] result_exp__77;
  wire is_result_nan__86;
  wire is_operand_inf__42;
  wire and_reduce_160339;
  wire [2:0] fraction_shift__404;
  wire [2:0] fraction_shift__301;
  wire is_subnormal__45;
  wire [7:0] high_exp__217;
  wire [7:0] result_exp__137;
  wire is_result_nan__125;
  wire is_operand_inf__61;
  wire and_reduce_160352;
  wire [2:0] fraction_shift__422;
  wire [2:0] fraction_shift__336;
  wire is_subnormal__65;
  wire [7:0] high_exp__286;
  wire [7:0] result_exp__197;
  wire [2:0] fraction_shift__369;
  wire [2:0] fraction_shift__232;
  wire [7:0] high_exp__89;
  wire [2:0] fraction_shift__33;
  wire result_sign__403;
  wire [7:0] result_exponent__11;
  wire result_sign__404;
  wire [2:0] fraction_shift__387;
  wire [2:0] fraction_shift__267;
  wire [7:0] high_exp__154;
  wire [2:0] fraction_shift__68;
  wire result_sign__500;
  wire [7:0] result_exponent__22;
  wire result_sign__501;
  wire [2:0] fraction_shift__405;
  wire [2:0] fraction_shift__302;
  wire [7:0] high_exp__218;
  wire [2:0] fraction_shift__125;
  wire result_sign__593;
  wire [7:0] result_exponent__41;
  wire result_sign__594;
  wire [2:0] fraction_shift__423;
  wire [2:0] fraction_shift__337;
  wire [7:0] high_exp__288;
  wire [2:0] fraction_shift__182;
  wire result_sign__699;
  wire [7:0] result_exponent__60;
  wire result_sign__700;
  wire [2:0] fraction_shift__6;
  wire result_sign__405;
  wire [7:0] result_exponent__1;
  wire [27:0] shrl_160412;
  wire [8:0] concat_160416;
  wire [2:0] fraction_shift__69;
  wire result_sign__502;
  wire [7:0] result_exponent__23;
  wire [27:0] shrl_160421;
  wire [8:0] concat_160425;
  wire [2:0] fraction_shift__126;
  wire result_sign__595;
  wire [7:0] result_exponent__42;
  wire [27:0] shrl_160430;
  wire [8:0] concat_160434;
  wire [2:0] fraction_shift__183;
  wire result_sign__701;
  wire [7:0] result_exponent__61;
  wire [27:0] shrl_160439;
  wire [8:0] concat_160443;
  wire [27:0] shrl_160444;
  wire [22:0] result_fraction__63;
  wire [22:0] result_fraction__66;
  wire [8:0] sum__11;
  wire [27:0] shrl_160452;
  wire [22:0] result_fraction__136;
  wire [22:0] result_fraction__142;
  wire [8:0] sum__24;
  wire [27:0] shrl_160460;
  wire [22:0] result_fraction__253;
  wire [22:0] result_fraction__259;
  wire [8:0] sum__43;
  wire [27:0] shrl_160468;
  wire [22:0] result_fraction__370;
  wire [22:0] result_fraction__376;
  wire [8:0] sum__62;
  wire [22:0] result_fraction__10;
  wire [8:0] sum__3;
  wire [22:0] result_fraction__64;
  wire [22:0] nan_fraction__83;
  wire [22:0] result_fraction__67;
  wire [22:0] nan_fraction__85;
  wire [22:0] result_fraction__137;
  wire [8:0] sum__25;
  wire [22:0] result_fraction__138;
  wire [22:0] nan_fraction__110;
  wire [22:0] result_fraction__144;
  wire [22:0] nan_fraction__112;
  wire [22:0] result_fraction__254;
  wire [8:0] sum__44;
  wire [22:0] result_fraction__255;
  wire [22:0] nan_fraction__137;
  wire [22:0] result_fraction__261;
  wire [22:0] nan_fraction__139;
  wire [22:0] result_fraction__371;
  wire [8:0] sum__63;
  wire [22:0] result_fraction__372;
  wire [22:0] nan_fraction__166;
  wire [22:0] result_fraction__378;
  wire [22:0] nan_fraction__168;
  wire [22:0] result_fraction__11;
  wire [22:0] nan_fraction__84;
  wire [22:0] result_fraction__65;
  wire [22:0] result_fraction__68;
  wire [7:0] prod_bexp__46;
  wire [7:0] x_bexp__692;
  wire [22:0] result_fraction__139;
  wire [22:0] nan_fraction__111;
  wire [22:0] result_fraction__140;
  wire [22:0] result_fraction__146;
  wire [7:0] prod_bexp__91;
  wire [7:0] x_bexp__693;
  wire [22:0] result_fraction__256;
  wire [22:0] nan_fraction__138;
  wire [22:0] result_fraction__257;
  wire [22:0] result_fraction__263;
  wire [7:0] prod_bexp__163;
  wire [7:0] x_bexp__694;
  wire [22:0] result_fraction__373;
  wire [22:0] nan_fraction__167;
  wire [22:0] result_fraction__374;
  wire [22:0] result_fraction__380;
  wire [7:0] prod_bexp__235;
  wire [7:0] x_bexp__695;
  wire [7:0] high_exp__351;
  wire [7:0] high_exp__352;
  wire [22:0] result_fraction__12;
  wire [7:0] prod_bexp__10;
  wire [7:0] x_bexp__696;
  wire fraction_is_zero__10;
  wire [22:0] prod_fraction__33;
  wire [7:0] incremented_sum__80;
  wire [7:0] high_exp__383;
  wire [7:0] high_exp__384;
  wire [22:0] result_fraction__141;
  wire [7:0] prod_bexp__92;
  wire [7:0] x_bexp__697;
  wire fraction_is_zero__22;
  wire [22:0] prod_fraction__67;
  wire [7:0] incremented_sum__98;
  wire [7:0] high_exp__415;
  wire [7:0] high_exp__416;
  wire [22:0] result_fraction__258;
  wire [7:0] prod_bexp__164;
  wire [7:0] x_bexp__698;
  wire fraction_is_zero__41;
  wire [22:0] prod_fraction__121;
  wire [7:0] incremented_sum__116;
  wire [7:0] high_exp__447;
  wire [7:0] high_exp__448;
  wire [22:0] result_fraction__375;
  wire [7:0] prod_bexp__236;
  wire [7:0] x_bexp__699;
  wire fraction_is_zero__60;
  wire [22:0] prod_fraction__175;
  wire [7:0] incremented_sum__134;
  wire fraction_is_zero__2;
  wire [22:0] prod_fraction__7;
  wire [7:0] incremented_sum__81;
  wire [27:0] wide_y__22;
  wire [7:0] x_bexpbs_difference__12;
  wire fraction_is_zero__23;
  wire [22:0] prod_fraction__68;
  wire [7:0] incremented_sum__99;
  wire [27:0] wide_y__47;
  wire [7:0] x_bexpbs_difference__23;
  wire fraction_is_zero__42;
  wire [22:0] prod_fraction__122;
  wire [7:0] incremented_sum__117;
  wire [27:0] wide_y__85;
  wire [7:0] x_bexpbs_difference__41;
  wire fraction_is_zero__61;
  wire [22:0] prod_fraction__176;
  wire [7:0] incremented_sum__135;
  wire [27:0] wide_y__123;
  wire [7:0] x_bexpbs_difference__59;
  wire [27:0] wide_y__5;
  wire [7:0] x_bexpbs_difference__3;
  wire [2:0] concat_160695;
  wire [7:0] x_bexp__94;
  wire [7:0] x_bexp__700;
  wire [27:0] wide_y__23;
  wire [7:0] sub_160701;
  wire [27:0] wide_y__48;
  wire [7:0] x_bexpbs_difference__24;
  wire [2:0] concat_160709;
  wire [7:0] x_bexp__187;
  wire [7:0] x_bexp__701;
  wire [27:0] wide_y__49;
  wire [7:0] sub_160715;
  wire [27:0] wide_y__86;
  wire [7:0] x_bexpbs_difference__42;
  wire [2:0] concat_160723;
  wire [7:0] x_bexp__331;
  wire [7:0] x_bexp__702;
  wire [27:0] wide_y__87;
  wire [7:0] sub_160729;
  wire [27:0] wide_y__124;
  wire [7:0] x_bexpbs_difference__60;
  wire [2:0] concat_160737;
  wire [7:0] x_bexp__475;
  wire [7:0] x_bexp__703;
  wire [27:0] wide_y__125;
  wire [7:0] sub_160743;
  wire [2:0] concat_160744;
  wire has_pos_inf__2;
  wire [7:0] x_bexp__22;
  wire [7:0] x_bexp__704;
  wire [27:0] wide_y__6;
  wire [7:0] sub_160751;
  wire result_sign__52;
  wire [22:0] x_fraction__94;
  wire [27:0] dropped__11;
  wire [2:0] concat_160759;
  wire has_pos_inf__23;
  wire [7:0] x_bexp__188;
  wire [7:0] x_bexp__705;
  wire [27:0] wide_y__50;
  wire [7:0] sub_160766;
  wire x_sign__45;
  wire result_sign__112;
  wire [22:0] x_fraction__187;
  wire [27:0] dropped__24;
  wire [2:0] concat_160775;
  wire has_pos_inf__42;
  wire [7:0] x_bexp__332;
  wire [7:0] x_bexp__706;
  wire [27:0] wide_y__88;
  wire [7:0] sub_160782;
  wire result_sign__209;
  wire [22:0] x_fraction__331;
  wire [27:0] dropped__43;
  wire [2:0] concat_160790;
  wire has_pos_inf__61;
  wire [7:0] x_bexp__476;
  wire [7:0] x_bexp__707;
  wire [27:0] wide_y__126;
  wire [7:0] sub_160797;
  wire x_sign__117;
  wire result_sign__306;
  wire [22:0] x_fraction__475;
  wire [27:0] dropped__62;
  wire result_sign__8;
  wire [22:0] x_fraction__22;
  wire [27:0] dropped__3;
  wire result_sign__53;
  wire [27:0] wide_x__22;
  wire result_sign__113;
  wire [22:0] x_fraction__188;
  wire [27:0] dropped__25;
  wire nand_160826;
  wire result_sign__118;
  wire result_sign__114;
  wire [27:0] wide_x__47;
  wire result_sign__210;
  wire [22:0] x_fraction__332;
  wire [27:0] dropped__44;
  wire result_sign__211;
  wire [27:0] wide_x__85;
  wire result_sign__307;
  wire [22:0] x_fraction__476;
  wire [27:0] dropped__63;
  wire nand_160854;
  wire result_sign__312;
  wire result_sign__308;
  wire [27:0] wide_x__123;
  wire result_sign__9;
  wire [27:0] wide_x__5;
  wire result_sign__54;
  wire [27:0] wide_x__23;
  wire result_sign__115;
  wire [27:0] wide_x__48;
  wire result_sign__120;
  wire result_sign__116;
  wire [27:0] wide_x__49;
  wire result_sign__212;
  wire [27:0] wide_x__86;
  wire result_sign__213;
  wire [27:0] wide_x__87;
  wire result_sign__309;
  wire [27:0] wide_x__124;
  wire result_sign__314;
  wire result_sign__310;
  wire [27:0] wide_x__125;
  wire result_sign__12;
  wire result_sign__10;
  wire [27:0] wide_x__6;
  wire x_sign__24;
  wire prod_sign__11;
  wire [27:0] neg_160911;
  wire [27:0] sticky__35;
  wire result_sign__121;
  wire result_sign__117;
  wire [27:0] wide_x__50;
  wire x_sign__47;
  wire prod_sign__23;
  wire [27:0] neg_160921;
  wire [27:0] sticky__76;
  wire result_sign__218;
  wire result_sign__214;
  wire [27:0] wide_x__88;
  wire x_sign__83;
  wire prod_sign__41;
  wire [27:0] neg_160931;
  wire [27:0] sticky__135;
  wire result_sign__315;
  wire result_sign__311;
  wire [27:0] wide_x__126;
  wire x_sign__119;
  wire prod_sign__59;
  wire [27:0] neg_160941;
  wire [27:0] sticky__194;
  wire x_sign__6;
  wire prod_sign__3;
  wire [27:0] neg_160946;
  wire [27:0] sticky__9;
  wire [27:0] xddend_y__11;
  wire x_sign__48;
  wire prod_sign__24;
  wire [27:0] neg_160955;
  wire [27:0] sticky__77;
  wire [27:0] xddend_y__23;
  wire x_sign__84;
  wire prod_sign__42;
  wire [27:0] neg_160964;
  wire [27:0] sticky__136;
  wire [27:0] xddend_y__41;
  wire x_sign__120;
  wire prod_sign__60;
  wire [27:0] neg_160973;
  wire [27:0] sticky__195;
  wire [27:0] xddend_y__59;
  wire [27:0] xddend_y__3;
  wire [24:0] sel_160984;
  wire result_sign__980;
  wire [27:0] xddend_y__24;
  wire [24:0] sel_160991;
  wire result_sign__981;
  wire [27:0] xddend_y__42;
  wire [24:0] sel_160998;
  wire result_sign__982;
  wire [27:0] xddend_y__60;
  wire [24:0] sel_161005;
  wire result_sign__983;
  wire [24:0] sel_161008;
  wire result_sign__984;
  wire [24:0] sel_161013;
  wire result_sign__985;
  wire [24:0] sel_161018;
  wire result_sign__986;
  wire [24:0] sel_161023;
  wire result_sign__987;
  wire [25:0] add_161030;
  wire [25:0] add_161033;
  wire [25:0] add_161036;
  wire [25:0] add_161039;
  wire [25:0] add_161040;
  wire [25:0] add_161043;
  wire [25:0] add_161046;
  wire [25:0] add_161049;
  wire [27:0] concat_161054;
  wire [27:0] concat_161057;
  wire [27:0] concat_161060;
  wire [27:0] concat_161063;
  wire [27:0] concat_161064;
  wire [27:0] concat_161067;
  wire [27:0] concat_161070;
  wire [27:0] concat_161073;
  wire [27:0] xbs_fraction__11;
  wire [27:0] xbs_fraction__23;
  wire [27:0] xbs_fraction__41;
  wire [27:0] xbs_fraction__59;
  wire [27:0] xbs_fraction__3;
  wire [27:0] reverse_161089;
  wire [27:0] xbs_fraction__24;
  wire [27:0] reverse_161091;
  wire [27:0] xbs_fraction__42;
  wire [27:0] reverse_161093;
  wire [27:0] xbs_fraction__60;
  wire [27:0] reverse_161095;
  wire [27:0] reverse_161096;
  wire [28:0] one_hot_161097;
  wire [27:0] reverse_161098;
  wire [28:0] one_hot_161099;
  wire [27:0] reverse_161100;
  wire [28:0] one_hot_161101;
  wire [27:0] reverse_161102;
  wire [28:0] one_hot_161103;
  wire [28:0] one_hot_161104;
  wire [4:0] encode_161105;
  wire [28:0] one_hot_161106;
  wire [4:0] encode_161107;
  wire [28:0] one_hot_161108;
  wire [4:0] encode_161109;
  wire [28:0] one_hot_161110;
  wire [4:0] encode_161111;
  wire [4:0] encode_161112;
  wire [4:0] encode_161114;
  wire [4:0] encode_161116;
  wire [4:0] encode_161118;
  wire cancel__12;
  wire carry_bit__11;
  wire [22:0] result_fraction__490;
  wire cancel__24;
  wire carry_bit__24;
  wire [22:0] result_fraction__557;
  wire cancel__43;
  wire carry_bit__43;
  wire [22:0] result_fraction__620;
  wire cancel__62;
  wire carry_bit__62;
  wire [22:0] result_fraction__691;
  wire cancel__3;
  wire carry_bit__3;
  wire [22:0] result_fraction__491;
  wire [27:0] leading_zeroes__11;
  wire cancel__25;
  wire carry_bit__25;
  wire [22:0] result_fraction__558;
  wire [27:0] leading_zeroes__24;
  wire cancel__44;
  wire carry_bit__44;
  wire [22:0] result_fraction__621;
  wire [27:0] leading_zeroes__43;
  wire cancel__63;
  wire carry_bit__63;
  wire [22:0] result_fraction__692;
  wire [27:0] leading_zeroes__62;
  wire [27:0] leading_zeroes__3;
  wire [26:0] carry_fraction__22;
  wire [27:0] add_161186;
  wire [27:0] leading_zeroes__25;
  wire [26:0] carry_fraction__47;
  wire [27:0] add_161199;
  wire [27:0] leading_zeroes__44;
  wire [31:0] array_index_161206;
  wire [26:0] carry_fraction__85;
  wire [27:0] add_161213;
  wire [27:0] leading_zeroes__63;
  wire [31:0] array_index_161220;
  wire [26:0] carry_fraction__123;
  wire [27:0] add_161227;
  wire [26:0] carry_fraction__5;
  wire [27:0] add_161234;
  wire [2:0] concat_161235;
  wire [26:0] carry_fraction__23;
  wire [26:0] cancel_fraction__11;
  wire [26:0] carry_fraction__48;
  wire [27:0] add_161244;
  wire [2:0] concat_161245;
  wire [26:0] carry_fraction__49;
  wire [26:0] cancel_fraction__24;
  wire [26:0] carry_fraction__86;
  wire [27:0] add_161254;
  wire [7:0] x_bexp__334;
  wire [2:0] concat_161256;
  wire [26:0] carry_fraction__87;
  wire [26:0] cancel_fraction__43;
  wire [26:0] carry_fraction__124;
  wire [27:0] add_161265;
  wire [7:0] x_bexp__478;
  wire [2:0] concat_161267;
  wire [26:0] carry_fraction__125;
  wire [26:0] cancel_fraction__62;
  wire [2:0] concat_161270;
  wire [26:0] carry_fraction__6;
  wire [26:0] cancel_fraction__3;
  wire result_sign__988;
  wire [26:0] shifted_fraction__11;
  wire [2:0] concat_161276;
  wire [26:0] carry_fraction__50;
  wire [26:0] cancel_fraction__25;
  wire [26:0] shifted_fraction__24;
  wire [2:0] concat_161280;
  wire [26:0] carry_fraction__88;
  wire [26:0] cancel_fraction__44;
  wire result_sign__989;
  wire [26:0] shifted_fraction__43;
  wire [2:0] concat_161286;
  wire [26:0] carry_fraction__126;
  wire [26:0] cancel_fraction__63;
  wire result_sign__990;
  wire [26:0] shifted_fraction__62;
  wire [26:0] shifted_fraction__3;
  wire result_sign__991;
  wire [26:0] shifted_fraction__25;
  wire result_sign__992;
  wire [26:0] shifted_fraction__44;
  wire result_sign__993;
  wire [26:0] shifted_fraction__63;
  wire result_sign__994;
  wire result_sign__995;
  wire result_sign__1105;
  wire [1:0] add_161313;
  wire [2:0] normal_chunk__11;
  wire [2:0] fraction_shift__233;
  wire [1:0] half_way_chunk__11;
  wire result_sign__996;
  wire [2:0] normal_chunk__24;
  wire [2:0] fraction_shift__268;
  wire [1:0] half_way_chunk__24;
  wire result_sign__997;
  wire result_sign__1109;
  wire [1:0] add_161332;
  wire [7:0] x_bexp__708;
  wire result_sign__598;
  wire [22:0] x_fraction__334;
  wire [2:0] normal_chunk__43;
  wire [2:0] fraction_shift__303;
  wire [1:0] half_way_chunk__43;
  wire result_sign__998;
  wire result_sign__1113;
  wire [1:0] add_161346;
  wire [7:0] x_bexp__709;
  wire result_sign__704;
  wire [22:0] x_fraction__478;
  wire [2:0] normal_chunk__62;
  wire [2:0] fraction_shift__338;
  wire [1:0] half_way_chunk__62;
  wire [2:0] normal_chunk__3;
  wire [2:0] fraction_shift__234;
  wire [1:0] half_way_chunk__3;
  wire result_sign__406;
  wire [24:0] add_161368;
  wire [2:0] normal_chunk__25;
  wire [2:0] fraction_shift__269;
  wire [1:0] half_way_chunk__25;
  wire result_sign__503;
  wire [24:0] add_161378;
  wire [2:0] normal_chunk__44;
  wire [2:0] fraction_shift__304;
  wire [1:0] half_way_chunk__44;
  wire ne_161387;
  wire result_sign__596;
  wire [24:0] add_161393;
  wire [2:0] normal_chunk__63;
  wire [2:0] fraction_shift__339;
  wire [1:0] half_way_chunk__63;
  wire ne_161402;
  wire result_sign__702;
  wire [24:0] add_161408;
  wire result_sign__407;
  wire [24:0] add_161412;
  wire [9:0] exp__13;
  wire do_round_up__23;
  wire result_sign__504;
  wire [24:0] add_161420;
  wire do_round_up__50;
  wire result_sign__597;
  wire [24:0] add_161427;
  wire [9:0] exp__190;
  wire [9:0] sign_ext_161429;
  wire [23:0] x_fraction__336;
  wire do_round_up__89;
  wire result_sign__703;
  wire [24:0] add_161438;
  wire [9:0] exp__272;
  wire [9:0] sign_ext_161440;
  wire [23:0] x_fraction__480;
  wire do_round_up__128;
  wire do_round_up__6;
  wire [9:0] exp__14;
  wire [27:0] rounded_fraction__11;
  wire do_round_up__51;
  wire [27:0] rounded_fraction__24;
  wire do_round_up__90;
  wire [9:0] exp__192;
  wire [23:0] x_fraction__338;
  wire result_sign__812;
  wire result_sign__813;
  wire [27:0] rounded_fraction__43;
  wire do_round_up__129;
  wire [9:0] exp__274;
  wire [23:0] x_fraction__482;
  wire result_sign__814;
  wire result_sign__815;
  wire [27:0] rounded_fraction__62;
  wire [27:0] rounded_fraction__3;
  wire result_sign__408;
  wire [7:0] x_bexp__578;
  wire rounding_carry__11;
  wire [27:0] rounded_fraction__25;
  wire result_sign__505;
  wire [7:0] x_bexp__596;
  wire rounding_carry__24;
  wire [27:0] rounded_fraction__44;
  wire [24:0] concat_161485;
  wire [24:0] concat_161486;
  wire result_sign__600;
  wire [7:0] x_bexp__614;
  wire rounding_carry__43;
  wire [27:0] rounded_fraction__63;
  wire [24:0] concat_161492;
  wire [24:0] concat_161493;
  wire result_sign__706;
  wire [7:0] x_bexp__632;
  wire rounding_carry__62;
  wire result_sign__409;
  wire [7:0] x_bexp__579;
  wire rounding_carry__3;
  wire [24:0] sel_161500;
  wire result_sign__506;
  wire [7:0] x_bexp__597;
  wire rounding_carry__25;
  wire result_sign__601;
  wire [7:0] x_bexp__615;
  wire rounding_carry__44;
  wire [24:0] sel_161511;
  wire result_sign__707;
  wire [7:0] x_bexp__633;
  wire rounding_carry__63;
  wire [24:0] sel_161517;
  wire result_sign__931;
  wire [22:0] fraction__33;
  wire result_sign__410;
  wire [8:0] add_161525;
  wire result_sign__507;
  wire [8:0] add_161531;
  wire result_sign__943;
  wire [22:0] fraction__424;
  wire result_sign__602;
  wire [8:0] add_161539;
  wire result_sign__951;
  wire [22:0] fraction__603;
  wire result_sign__708;
  wire [8:0] add_161547;
  wire result_sign__411;
  wire [8:0] add_161551;
  wire [23:0] fraction__34;
  wire result_sign__508;
  wire [8:0] add_161564;
  wire result_sign__603;
  wire [8:0] add_161573;
  wire [23:0] fraction__426;
  wire result_sign__709;
  wire [8:0] add_161586;
  wire [23:0] fraction__605;
  wire do_round_up__7;
  wire [23:0] add_161604;
  wire [9:0] add_161605;
  wire [9:0] add_161613;
  wire do_round_up__92;
  wire [23:0] add_161622;
  wire [9:0] add_161623;
  wire do_round_up__131;
  wire [23:0] add_161632;
  wire [9:0] add_161633;
  wire [9:0] add_161636;
  wire [23:0] fraction__35;
  wire [9:0] wide_exponent__33;
  wire [9:0] add_161643;
  wire [9:0] wide_exponent__70;
  wire [9:0] add_161648;
  wire [23:0] fraction__428;
  wire [9:0] wide_exponent__127;
  wire [9:0] add_161655;
  wire [23:0] fraction__607;
  wire [9:0] wide_exponent__184;
  wire [9:0] wide_exponent__7;
  wire [9:0] add_161665;
  wire [9:0] wide_exponent__34;
  wire [9:0] wide_exponent__71;
  wire [9:0] wide_exponent__72;
  wire [9:0] wide_exponent__128;
  wire [9:0] add_161673;
  wire [9:0] wide_exponent__129;
  wire [9:0] wide_exponent__185;
  wire [9:0] add_161678;
  wire [9:0] wide_exponent__186;
  wire [9:0] wide_exponent__8;
  wire [9:0] exp__16;
  wire [7:0] high_exp__367;
  wire [22:0] result_fraction__773;
  wire [7:0] high_exp__368;
  wire [22:0] result_fraction__774;
  wire [7:0] high_exp__91;
  wire [22:0] result_fraction__492;
  wire [7:0] high_exp__92;
  wire [22:0] result_fraction__493;
  wire [9:0] wide_exponent__73;
  wire [7:0] high_exp__399;
  wire [22:0] result_fraction__806;
  wire [7:0] high_exp__400;
  wire [22:0] result_fraction__807;
  wire [7:0] high_exp__156;
  wire [22:0] result_fraction__559;
  wire [7:0] high_exp__157;
  wire [22:0] result_fraction__560;
  wire [9:0] wide_exponent__130;
  wire [9:0] exp__196;
  wire [7:0] high_exp__431;
  wire [22:0] result_fraction__839;
  wire [7:0] high_exp__432;
  wire [22:0] result_fraction__840;
  wire [7:0] high_exp__220;
  wire [22:0] result_fraction__622;
  wire [7:0] high_exp__221;
  wire [22:0] result_fraction__623;
  wire [9:0] wide_exponent__187;
  wire [9:0] exp__278;
  wire [7:0] high_exp__463;
  wire [22:0] result_fraction__872;
  wire [7:0] high_exp__464;
  wire [22:0] result_fraction__873;
  wire [7:0] high_exp__290;
  wire [22:0] result_fraction__693;
  wire [7:0] high_exp__291;
  wire [22:0] result_fraction__694;
  wire [7:0] high_exp__353;
  wire [22:0] result_fraction__758;
  wire [7:0] high_exp__354;
  wire [22:0] result_fraction__759;
  wire [7:0] high_exp__93;
  wire [22:0] result_fraction__494;
  wire [7:0] high_exp__94;
  wire [22:0] result_fraction__495;
  wire ne_161738;
  wire ne_161740;
  wire eq_161741;
  wire eq_161742;
  wire eq_161743;
  wire eq_161744;
  wire [7:0] high_exp__385;
  wire [22:0] result_fraction__791;
  wire [7:0] high_exp__386;
  wire [22:0] result_fraction__792;
  wire [7:0] high_exp__158;
  wire [22:0] result_fraction__561;
  wire [7:0] high_exp__159;
  wire [22:0] result_fraction__562;
  wire ne_161756;
  wire ne_161758;
  wire eq_161759;
  wire eq_161760;
  wire eq_161761;
  wire eq_161762;
  wire [7:0] high_exp__417;
  wire [22:0] result_fraction__824;
  wire [7:0] high_exp__418;
  wire [22:0] result_fraction__825;
  wire [7:0] high_exp__222;
  wire [22:0] result_fraction__624;
  wire [7:0] high_exp__223;
  wire [22:0] result_fraction__625;
  wire ne_161775;
  wire ne_161777;
  wire eq_161778;
  wire eq_161779;
  wire eq_161780;
  wire eq_161781;
  wire [7:0] high_exp__449;
  wire [22:0] result_fraction__857;
  wire [7:0] high_exp__450;
  wire [22:0] result_fraction__858;
  wire [7:0] high_exp__292;
  wire [22:0] result_fraction__695;
  wire [7:0] high_exp__293;
  wire [22:0] result_fraction__696;
  wire ne_161794;
  wire ne_161796;
  wire eq_161797;
  wire eq_161798;
  wire eq_161799;
  wire eq_161800;
  wire ne_161803;
  wire ne_161805;
  wire eq_161806;
  wire eq_161807;
  wire eq_161808;
  wire eq_161809;
  wire [8:0] result_exp__10;
  wire ne_161820;
  wire ne_161822;
  wire eq_161823;
  wire eq_161824;
  wire eq_161825;
  wire eq_161826;
  wire ne_161835;
  wire ne_161837;
  wire eq_161838;
  wire eq_161839;
  wire eq_161840;
  wire eq_161841;
  wire [8:0] result_exp__140;
  wire ne_161852;
  wire ne_161854;
  wire eq_161855;
  wire eq_161856;
  wire eq_161857;
  wire eq_161858;
  wire [8:0] result_exp__200;
  wire [8:0] result_exp__11;
  wire [8:0] wide_exponent__35;
  wire has_pos_inf__11;
  wire has_neg_inf__11;
  wire [8:0] wide_exponent__74;
  wire has_pos_inf__24;
  wire has_neg_inf__24;
  wire [7:0] high_exp__226;
  wire [22:0] result_fraction__627;
  wire [22:0] result_fraction__626;
  wire [8:0] result_exp__142;
  wire [8:0] wide_exponent__131;
  wire has_pos_inf__43;
  wire has_neg_inf__43;
  wire [7:0] high_exp__296;
  wire [22:0] result_fraction__698;
  wire [22:0] result_fraction__697;
  wire [8:0] result_exp__202;
  wire [8:0] wide_exponent__188;
  wire has_pos_inf__62;
  wire has_neg_inf__62;
  wire [8:0] wide_exponent__9;
  wire has_pos_inf__3;
  wire has_neg_inf__3;
  wire [8:0] wide_exponent__75;
  wire has_pos_inf__25;
  wire has_neg_inf__25;
  wire [8:0] wide_exponent__132;
  wire has_pos_inf__44;
  wire has_neg_inf__44;
  wire is_result_nan__91;
  wire ne_161937;
  wire [8:0] wide_exponent__189;
  wire has_pos_inf__63;
  wire has_neg_inf__63;
  wire is_result_nan__130;
  wire ne_161951;
  wire and_reduce_161969;
  wire is_result_nan__23;
  wire is_operand_inf__11;
  wire and_reduce_161975;
  wire is_result_nan__50;
  wire is_operand_inf__24;
  wire and_reduce_161988;
  wire is_result_nan__92;
  wire has_inf_arg__47;
  wire and_reduce_161999;
  wire is_result_nan__89;
  wire is_operand_inf__43;
  wire and_reduce_162005;
  wire is_result_nan__131;
  wire has_inf_arg__67;
  wire and_reduce_162016;
  wire is_result_nan__128;
  wire is_operand_inf__62;
  wire and_reduce_162022;
  wire is_result_nan__6;
  wire is_operand_inf__3;
  wire and_reduce_162029;
  wire [7:0] high_exp__97;
  wire [2:0] fraction_shift__370;
  wire [2:0] fraction_shift__235;
  wire [7:0] high_exp__95;
  wire [7:0] result_exp__38;
  wire is_result_nan__51;
  wire is_operand_inf__25;
  wire and_reduce_162043;
  wire [2:0] fraction_shift__388;
  wire [2:0] fraction_shift__270;
  wire [7:0] high_exp__160;
  wire is_result_nan__90;
  wire is_operand_inf__44;
  wire and_reduce_162055;
  wire [7:0] high_exp__227;
  wire [2:0] fraction_shift__406;
  wire [2:0] fraction_shift__305;
  wire [7:0] high_exp__224;
  wire [7:0] result_exp__143;
  wire is_result_nan__129;
  wire is_operand_inf__63;
  wire and_reduce_162070;
  wire [7:0] high_exp__297;
  wire [2:0] fraction_shift__424;
  wire [2:0] fraction_shift__340;
  wire [7:0] high_exp__294;
  wire [7:0] result_exp__203;
  wire [2:0] fraction_shift__371;
  wire [2:0] fraction_shift__236;
  wire is_subnormal__4;
  wire [7:0] high_exp__96;
  wire [7:0] result_exp__12;
  wire [2:0] fraction_shift__36;
  wire result_sign__412;
  wire [7:0] result_exponent__12;
  wire result_sign__413;
  wire [2:0] fraction_shift__389;
  wire [2:0] fraction_shift__271;
  wire [7:0] high_exp__161;
  wire [2:0] fraction_shift__74;
  wire result_sign__509;
  wire [7:0] result_exponent__24;
  wire [2:0] fraction_shift__407;
  wire [2:0] fraction_shift__306;
  wire is_subnormal__48;
  wire [7:0] high_exp__225;
  wire [7:0] result_exp__144;
  wire [2:0] fraction_shift__131;
  wire result_sign__604;
  wire [7:0] result_exponent__43;
  wire result_sign__605;
  wire [2:0] fraction_shift__425;
  wire [2:0] fraction_shift__341;
  wire is_subnormal__68;
  wire [7:0] high_exp__295;
  wire [7:0] result_exp__204;
  wire [2:0] fraction_shift__188;
  wire result_sign__710;
  wire [7:0] result_exponent__62;
  wire result_sign__711;
  wire [2:0] fraction_shift__9;
  wire result_sign__414;
  wire [7:0] result_exponent__3;
  wire result_sign__415;
  wire [27:0] shrl_162134;
  wire [2:0] fraction_shift__75;
  wire result_sign__510;
  wire [7:0] result_exponent__25;
  wire [27:0] shrl_162142;
  wire [2:0] fraction_shift__132;
  wire result_sign__606;
  wire [7:0] result_exponent__44;
  wire result_sign__607;
  wire [27:0] shrl_162152;
  wire [2:0] fraction_shift__189;
  wire result_sign__712;
  wire [7:0] result_exponent__63;
  wire result_sign__713;
  wire [27:0] shrl_162163;
  wire [8:0] concat_162166;
  wire [27:0] shrl_162167;
  wire [22:0] result_fraction__69;
  wire [8:0] sum__12;
  wire [27:0] shrl_162175;
  wire [22:0] result_fraction__148;
  wire [8:0] sum__26;
  wire [27:0] shrl_162181;
  wire [22:0] result_fraction__265;
  wire [8:0] sum__45;
  wire [27:0] shrl_162189;
  wire [8:0] concat_162193;
  wire [22:0] result_fraction__382;
  wire [8:0] sum__64;
  wire [22:0] result_fraction__16;
  wire [22:0] result_fraction__19;
  wire [8:0] sum__4;
  wire [22:0] result_fraction__70;
  wire [22:0] nan_fraction__86;
  wire [22:0] result_fraction__149;
  wire [8:0] sum__27;
  wire [22:0] result_fraction__150;
  wire [22:0] nan_fraction__113;
  wire [22:0] result_fraction__266;
  wire [22:0] result_fraction__272;
  wire [8:0] sum__46;
  wire [22:0] result_fraction__267;
  wire [22:0] nan_fraction__140;
  wire [22:0] result_fraction__383;
  wire [22:0] result_fraction__389;
  wire [8:0] sum__65;
  wire [22:0] result_fraction__384;
  wire [22:0] nan_fraction__169;
  wire [22:0] result_fraction__17;
  wire [22:0] nan_fraction__87;
  wire [22:0] result_fraction__20;
  wire [22:0] nan_fraction__88;
  wire [22:0] result_fraction__71;
  wire [22:0] result_fraction__473;
  wire [7:0] prod_bexp__50;
  wire [7:0] x_bexp__710;
  wire [22:0] result_fraction__151;
  wire [22:0] nan_fraction__114;
  wire [22:0] result_fraction__152;
  wire [7:0] prod_bexp__99;
  wire [7:0] x_bexp__711;
  wire [22:0] result_fraction__268;
  wire [22:0] nan_fraction__141;
  wire [22:0] result_fraction__274;
  wire [22:0] nan_fraction__142;
  wire [22:0] result_fraction__269;
  wire [22:0] result_fraction__474;
  wire [7:0] prod_bexp__171;
  wire [7:0] x_bexp__712;
  wire [22:0] result_fraction__385;
  wire [22:0] nan_fraction__170;
  wire [22:0] result_fraction__391;
  wire [22:0] nan_fraction__171;
  wire [22:0] result_fraction__386;
  wire [22:0] result_fraction__475;
  wire [7:0] prod_bexp__243;
  wire [7:0] x_bexp__713;
  wire [22:0] result_fraction__18;
  wire [22:0] result_fraction__21;
  wire [7:0] prod_bexp__14;
  wire [7:0] x_bexp__714;
  wire fraction_is_zero__11;
  wire [22:0] prod_fraction__36;
  wire [7:0] incremented_sum__82;
  wire [22:0] result_fraction__153;
  wire [7:0] prod_bexp__100;
  wire [7:0] x_bexp__715;
  wire fraction_is_zero__24;
  wire [22:0] prod_fraction__73;
  wire [7:0] incremented_sum__100;
  wire [22:0] result_fraction__270;
  wire [22:0] result_fraction__276;
  wire [7:0] prod_bexp__172;
  wire [7:0] x_bexp__716;
  wire fraction_is_zero__43;
  wire [22:0] prod_fraction__127;
  wire [7:0] incremented_sum__118;
  wire [22:0] result_fraction__387;
  wire [22:0] result_fraction__393;
  wire [7:0] prod_bexp__244;
  wire [7:0] x_bexp__717;
  wire fraction_is_zero__62;
  wire [22:0] prod_fraction__181;
  wire [7:0] incremented_sum__136;
  wire fraction_is_zero__3;
  wire [22:0] prod_fraction__10;
  wire [7:0] incremented_sum__83;
  wire [27:0] wide_y__24;
  wire [7:0] x_bexpbs_difference__13;
  wire fraction_is_zero__25;
  wire [22:0] prod_fraction__74;
  wire [7:0] incremented_sum__101;
  wire [27:0] wide_y__51;
  wire [7:0] x_bexpbs_difference__25;
  wire fraction_is_zero__44;
  wire [22:0] prod_fraction__128;
  wire [7:0] incremented_sum__119;
  wire [27:0] wide_y__89;
  wire [7:0] x_bexpbs_difference__43;
  wire fraction_is_zero__63;
  wire [22:0] prod_fraction__182;
  wire [7:0] incremented_sum__137;
  wire [27:0] wide_y__127;
  wire [7:0] x_bexpbs_difference__61;
  wire [27:0] wide_y__7;
  wire [7:0] x_bexpbs_difference__4;
  wire [2:0] concat_162407;
  wire [7:0] x_bexp__102;
  wire [7:0] x_bexp__718;
  wire [27:0] wide_y__25;
  wire [7:0] sub_162413;
  wire [27:0] wide_y__52;
  wire [7:0] x_bexpbs_difference__26;
  wire [2:0] concat_162419;
  wire [7:0] x_bexp__203;
  wire [7:0] x_bexp__719;
  wire [27:0] wide_y__53;
  wire [7:0] sub_162425;
  wire [27:0] wide_y__90;
  wire [7:0] x_bexpbs_difference__44;
  wire [2:0] concat_162431;
  wire [7:0] x_bexp__347;
  wire [7:0] x_bexp__720;
  wire [27:0] wide_y__91;
  wire [7:0] sub_162437;
  wire [27:0] wide_y__128;
  wire [7:0] x_bexpbs_difference__62;
  wire [2:0] concat_162443;
  wire [7:0] x_bexp__491;
  wire [7:0] x_bexp__721;
  wire [27:0] wide_y__129;
  wire [7:0] sub_162449;
  wire [2:0] concat_162450;
  wire [7:0] x_bexp__30;
  wire [7:0] x_bexp__722;
  wire [27:0] wide_y__8;
  wire [7:0] sub_162456;
  wire [7:0] high_exp__480;
  wire result_sign__57;
  wire [22:0] x_fraction__102;
  wire [27:0] dropped__12;
  wire [2:0] concat_162465;
  wire [7:0] x_bexp__204;
  wire [7:0] x_bexp__723;
  wire [27:0] wide_y__54;
  wire [7:0] sub_162471;
  wire result_sign__122;
  wire [22:0] x_fraction__203;
  wire [27:0] dropped__26;
  wire [2:0] concat_162479;
  wire [7:0] x_bexp__348;
  wire [7:0] x_bexp__724;
  wire [27:0] wide_y__92;
  wire [7:0] sub_162485;
  wire [7:0] high_exp__484;
  wire result_sign__219;
  wire [22:0] x_fraction__347;
  wire [27:0] dropped__45;
  wire [2:0] concat_162494;
  wire [7:0] x_bexp__492;
  wire [7:0] x_bexp__725;
  wire [27:0] wide_y__130;
  wire [7:0] sub_162500;
  wire [7:0] high_exp__487;
  wire result_sign__316;
  wire [22:0] x_fraction__491;
  wire [27:0] dropped__64;
  wire result_sign__13;
  wire [22:0] x_fraction__30;
  wire [27:0] dropped__4;
  wire result_sign__58;
  wire [27:0] wide_x__24;
  wire result_sign__123;
  wire [22:0] x_fraction__204;
  wire [27:0] dropped__27;
  wire result_sign__124;
  wire [27:0] wide_x__51;
  wire x_sign__86;
  wire result_sign__220;
  wire [22:0] x_fraction__348;
  wire [27:0] dropped__46;
  wire result_sign__221;
  wire [27:0] wide_x__89;
  wire x_sign__122;
  wire result_sign__317;
  wire [22:0] x_fraction__492;
  wire [27:0] dropped__65;
  wire result_sign__318;
  wire [27:0] wide_x__127;
  wire result_sign__14;
  wire [27:0] wide_x__7;
  wire result_sign__61;
  wire result_sign__59;
  wire [27:0] wide_x__25;
  wire result_sign__125;
  wire [27:0] wide_x__52;
  wire result_sign__126;
  wire [27:0] wide_x__53;
  wire nand_162587;
  wire result_sign__226;
  wire result_sign__222;
  wire [27:0] wide_x__90;
  wire result_sign__227;
  wire result_sign__223;
  wire [27:0] wide_x__91;
  wire nand_162600;
  wire result_sign__323;
  wire result_sign__319;
  wire [27:0] wide_x__128;
  wire result_sign__324;
  wire result_sign__320;
  wire [27:0] wide_x__129;
  wire result_sign__15;
  wire [27:0] wide_x__8;
  wire x_sign__26;
  wire prod_sign__12;
  wire [27:0] neg_162619;
  wire [27:0] sticky__38;
  wire result_sign__127;
  wire [27:0] wide_x__54;
  wire x_sign__51;
  wire prod_sign__25;
  wire [27:0] neg_162628;
  wire [27:0] sticky__82;
  wire result_sign__228;
  wire result_sign__224;
  wire [27:0] wide_x__92;
  wire x_sign__87;
  wire prod_sign__43;
  wire [27:0] neg_162638;
  wire [27:0] sticky__141;
  wire result_sign__325;
  wire result_sign__321;
  wire [27:0] wide_x__130;
  wire x_sign__123;
  wire prod_sign__61;
  wire [27:0] neg_162648;
  wire [27:0] sticky__200;
  wire x_sign__8;
  wire prod_sign__4;
  wire [27:0] neg_162653;
  wire [27:0] sticky__12;
  wire [27:0] xddend_y__12;
  wire x_sign__52;
  wire prod_sign__26;
  wire [27:0] neg_162662;
  wire [27:0] sticky__83;
  wire [27:0] xddend_y__25;
  wire x_sign__88;
  wire prod_sign__44;
  wire [27:0] neg_162671;
  wire [27:0] sticky__142;
  wire [27:0] xddend_y__43;
  wire x_sign__124;
  wire prod_sign__62;
  wire [27:0] neg_162680;
  wire [27:0] sticky__201;
  wire [27:0] xddend_y__61;
  wire [27:0] xddend_y__4;
  wire [24:0] sel_162691;
  wire result_sign__999;
  wire [27:0] xddend_y__26;
  wire [24:0] sel_162698;
  wire result_sign__1000;
  wire [27:0] xddend_y__44;
  wire [24:0] sel_162705;
  wire result_sign__1001;
  wire [27:0] xddend_y__62;
  wire [24:0] sel_162712;
  wire result_sign__1002;
  wire [24:0] sel_162715;
  wire result_sign__1003;
  wire [24:0] sel_162720;
  wire result_sign__1004;
  wire [24:0] sel_162725;
  wire result_sign__1005;
  wire [24:0] sel_162730;
  wire result_sign__1006;
  wire [25:0] add_162737;
  wire [25:0] add_162740;
  wire [25:0] add_162743;
  wire [25:0] add_162746;
  wire [25:0] add_162747;
  wire [25:0] add_162750;
  wire [25:0] add_162753;
  wire [25:0] add_162756;
  wire [27:0] concat_162761;
  wire [27:0] concat_162764;
  wire [27:0] concat_162767;
  wire [27:0] concat_162770;
  wire [27:0] concat_162771;
  wire [27:0] concat_162774;
  wire [27:0] concat_162777;
  wire [27:0] concat_162780;
  wire [27:0] xbs_fraction__12;
  wire [27:0] xbs_fraction__25;
  wire [27:0] xbs_fraction__43;
  wire [27:0] xbs_fraction__61;
  wire [27:0] xbs_fraction__4;
  wire [27:0] reverse_162796;
  wire [27:0] xbs_fraction__26;
  wire [27:0] reverse_162798;
  wire [27:0] xbs_fraction__44;
  wire [27:0] reverse_162800;
  wire [27:0] xbs_fraction__62;
  wire [27:0] reverse_162802;
  wire [27:0] reverse_162803;
  wire [28:0] one_hot_162804;
  wire [27:0] reverse_162805;
  wire [28:0] one_hot_162806;
  wire [27:0] reverse_162807;
  wire [28:0] one_hot_162808;
  wire [27:0] reverse_162809;
  wire [28:0] one_hot_162810;
  wire [28:0] one_hot_162811;
  wire [4:0] encode_162812;
  wire [28:0] one_hot_162813;
  wire [4:0] encode_162814;
  wire [28:0] one_hot_162815;
  wire [4:0] encode_162816;
  wire [28:0] one_hot_162817;
  wire [4:0] encode_162818;
  wire [4:0] encode_162819;
  wire [4:0] encode_162821;
  wire [4:0] encode_162823;
  wire [4:0] encode_162825;
  wire cancel__13;
  wire carry_bit__12;
  wire [22:0] result_fraction__496;
  wire cancel__26;
  wire carry_bit__26;
  wire [22:0] result_fraction__563;
  wire cancel__45;
  wire carry_bit__45;
  wire [22:0] result_fraction__628;
  wire cancel__64;
  wire carry_bit__64;
  wire [22:0] result_fraction__699;
  wire cancel__4;
  wire carry_bit__4;
  wire [22:0] result_fraction__497;
  wire [27:0] leading_zeroes__12;
  wire cancel__27;
  wire carry_bit__27;
  wire [22:0] result_fraction__564;
  wire [27:0] leading_zeroes__26;
  wire cancel__46;
  wire carry_bit__46;
  wire [22:0] result_fraction__629;
  wire [27:0] leading_zeroes__45;
  wire cancel__65;
  wire carry_bit__65;
  wire [22:0] result_fraction__700;
  wire [27:0] leading_zeroes__64;
  wire [27:0] leading_zeroes__4;
  wire [26:0] carry_fraction__24;
  wire [27:0] add_162891;
  wire [27:0] leading_zeroes__27;
  wire [26:0] carry_fraction__51;
  wire [27:0] add_162904;
  wire [27:0] leading_zeroes__46;
  wire [26:0] carry_fraction__89;
  wire [27:0] add_162917;
  wire [27:0] leading_zeroes__65;
  wire [26:0] carry_fraction__127;
  wire [27:0] add_162930;
  wire [26:0] carry_fraction__7;
  wire [27:0] add_162937;
  wire [2:0] concat_162938;
  wire [26:0] carry_fraction__25;
  wire [26:0] cancel_fraction__12;
  wire [26:0] carry_fraction__52;
  wire [27:0] add_162947;
  wire [2:0] concat_162948;
  wire [26:0] carry_fraction__53;
  wire [26:0] cancel_fraction__26;
  wire [26:0] carry_fraction__90;
  wire [27:0] add_162957;
  wire [2:0] concat_162958;
  wire [26:0] carry_fraction__91;
  wire [26:0] cancel_fraction__45;
  wire [26:0] carry_fraction__128;
  wire [27:0] add_162967;
  wire [2:0] concat_162968;
  wire [26:0] carry_fraction__129;
  wire [26:0] cancel_fraction__64;
  wire [2:0] concat_162971;
  wire [26:0] carry_fraction__8;
  wire [26:0] cancel_fraction__4;
  wire [26:0] shifted_fraction__12;
  wire [2:0] concat_162975;
  wire [26:0] carry_fraction__54;
  wire [26:0] cancel_fraction__27;
  wire [26:0] shifted_fraction__26;
  wire [2:0] concat_162979;
  wire [26:0] carry_fraction__92;
  wire [26:0] cancel_fraction__46;
  wire [26:0] shifted_fraction__45;
  wire [2:0] concat_162983;
  wire [26:0] carry_fraction__130;
  wire [26:0] cancel_fraction__65;
  wire [26:0] shifted_fraction__64;
  wire [26:0] shifted_fraction__4;
  wire result_sign__1007;
  wire [26:0] shifted_fraction__27;
  wire result_sign__1008;
  wire [26:0] shifted_fraction__46;
  wire result_sign__1009;
  wire [26:0] shifted_fraction__65;
  wire result_sign__1010;
  wire result_sign__1011;
  wire [2:0] normal_chunk__12;
  wire [2:0] fraction_shift__237;
  wire [1:0] half_way_chunk__12;
  wire result_sign__1012;
  wire [2:0] normal_chunk__26;
  wire [2:0] fraction_shift__272;
  wire [1:0] half_way_chunk__26;
  wire result_sign__1013;
  wire [2:0] normal_chunk__45;
  wire [2:0] fraction_shift__307;
  wire [1:0] half_way_chunk__45;
  wire result_sign__1014;
  wire [2:0] normal_chunk__64;
  wire [2:0] fraction_shift__342;
  wire [1:0] half_way_chunk__64;
  wire [2:0] normal_chunk__4;
  wire [2:0] fraction_shift__238;
  wire [1:0] half_way_chunk__4;
  wire result_sign__416;
  wire [24:0] add_163040;
  wire [2:0] normal_chunk__27;
  wire [2:0] fraction_shift__273;
  wire [1:0] half_way_chunk__27;
  wire result_sign__511;
  wire [24:0] add_163050;
  wire [2:0] normal_chunk__46;
  wire [2:0] fraction_shift__308;
  wire [1:0] half_way_chunk__46;
  wire result_sign__608;
  wire [24:0] add_163060;
  wire [2:0] normal_chunk__65;
  wire [2:0] fraction_shift__343;
  wire [1:0] half_way_chunk__65;
  wire result_sign__714;
  wire [24:0] add_163070;
  wire result_sign__417;
  wire [24:0] add_163074;
  wire do_round_up__25;
  wire result_sign__512;
  wire [24:0] add_163081;
  wire do_round_up__54;
  wire result_sign__609;
  wire [24:0] add_163088;
  wire do_round_up__93;
  wire result_sign__715;
  wire [24:0] add_163095;
  wire do_round_up__132;
  wire do_round_up__8;
  wire [27:0] rounded_fraction__12;
  wire do_round_up__55;
  wire [27:0] rounded_fraction__26;
  wire do_round_up__94;
  wire [27:0] rounded_fraction__45;
  wire do_round_up__133;
  wire [27:0] rounded_fraction__64;
  wire [27:0] rounded_fraction__4;
  wire result_sign__418;
  wire [7:0] x_bexp__580;
  wire rounding_carry__12;
  wire [27:0] rounded_fraction__27;
  wire result_sign__513;
  wire [7:0] x_bexp__598;
  wire rounding_carry__26;
  wire [27:0] rounded_fraction__46;
  wire result_sign__610;
  wire [7:0] x_bexp__616;
  wire rounding_carry__45;
  wire [27:0] rounded_fraction__65;
  wire result_sign__716;
  wire [7:0] x_bexp__634;
  wire rounding_carry__64;
  wire result_sign__419;
  wire [7:0] x_bexp__581;
  wire rounding_carry__4;
  wire result_sign__514;
  wire [7:0] x_bexp__599;
  wire rounding_carry__27;
  wire result_sign__611;
  wire [7:0] x_bexp__617;
  wire rounding_carry__46;
  wire result_sign__717;
  wire [7:0] x_bexp__635;
  wire rounding_carry__65;
  wire result_sign__420;
  wire [8:0] add_163154;
  wire result_sign__515;
  wire [8:0] add_163160;
  wire result_sign__612;
  wire [8:0] add_163166;
  wire result_sign__718;
  wire [8:0] add_163172;
  wire result_sign__421;
  wire [8:0] add_163176;
  wire result_sign__516;
  wire [8:0] add_163185;
  wire result_sign__613;
  wire [8:0] add_163194;
  wire result_sign__719;
  wire [8:0] add_163203;
  wire [9:0] add_163216;
  wire [9:0] add_163224;
  wire [9:0] add_163232;
  wire [9:0] add_163240;
  wire [9:0] add_163243;
  wire [9:0] wide_exponent__36;
  wire [9:0] add_163248;
  wire [9:0] wide_exponent__76;
  wire [9:0] add_163253;
  wire [9:0] wide_exponent__133;
  wire [9:0] add_163258;
  wire [9:0] wide_exponent__190;
  wire [9:0] wide_exponent__10;
  wire [9:0] wide_exponent__37;
  wire [9:0] wide_exponent__77;
  wire [9:0] wide_exponent__78;
  wire [9:0] wide_exponent__134;
  wire [9:0] wide_exponent__135;
  wire [9:0] wide_exponent__191;
  wire [9:0] wide_exponent__192;
  wire [9:0] wide_exponent__11;
  wire [7:0] high_exp__369;
  wire [22:0] result_fraction__775;
  wire [7:0] high_exp__370;
  wire [22:0] result_fraction__776;
  wire [7:0] high_exp__98;
  wire [22:0] result_fraction__498;
  wire [7:0] high_exp__99;
  wire [22:0] result_fraction__499;
  wire [9:0] wide_exponent__79;
  wire [7:0] high_exp__401;
  wire [22:0] result_fraction__808;
  wire [7:0] high_exp__402;
  wire [22:0] result_fraction__809;
  wire [7:0] high_exp__162;
  wire [22:0] result_fraction__565;
  wire [7:0] high_exp__163;
  wire [22:0] result_fraction__566;
  wire [9:0] wide_exponent__136;
  wire [7:0] high_exp__433;
  wire [22:0] result_fraction__841;
  wire [7:0] high_exp__434;
  wire [22:0] result_fraction__842;
  wire [7:0] high_exp__228;
  wire [22:0] result_fraction__630;
  wire [7:0] high_exp__229;
  wire [22:0] result_fraction__631;
  wire [9:0] wide_exponent__193;
  wire [7:0] high_exp__465;
  wire [22:0] result_fraction__874;
  wire [7:0] high_exp__466;
  wire [22:0] result_fraction__875;
  wire [7:0] high_exp__298;
  wire [22:0] result_fraction__701;
  wire [7:0] high_exp__299;
  wire [22:0] result_fraction__702;
  wire [7:0] high_exp__355;
  wire [22:0] result_fraction__760;
  wire [7:0] high_exp__356;
  wire [22:0] result_fraction__761;
  wire [7:0] high_exp__100;
  wire [22:0] result_fraction__500;
  wire [7:0] high_exp__101;
  wire [22:0] result_fraction__501;
  wire ne_163326;
  wire ne_163328;
  wire eq_163329;
  wire eq_163330;
  wire eq_163331;
  wire eq_163332;
  wire [7:0] high_exp__387;
  wire [22:0] result_fraction__793;
  wire [7:0] high_exp__388;
  wire [22:0] result_fraction__794;
  wire [7:0] high_exp__164;
  wire [22:0] result_fraction__567;
  wire [7:0] high_exp__165;
  wire [22:0] result_fraction__568;
  wire ne_163344;
  wire ne_163346;
  wire eq_163347;
  wire eq_163348;
  wire eq_163349;
  wire eq_163350;
  wire [7:0] high_exp__419;
  wire [22:0] result_fraction__826;
  wire [7:0] high_exp__420;
  wire [22:0] result_fraction__827;
  wire [7:0] high_exp__230;
  wire [22:0] result_fraction__632;
  wire [7:0] high_exp__231;
  wire [22:0] result_fraction__633;
  wire ne_163362;
  wire ne_163364;
  wire eq_163365;
  wire eq_163366;
  wire eq_163367;
  wire eq_163368;
  wire [7:0] high_exp__451;
  wire [22:0] result_fraction__859;
  wire [7:0] high_exp__452;
  wire [22:0] result_fraction__860;
  wire [7:0] high_exp__300;
  wire [22:0] result_fraction__703;
  wire [7:0] high_exp__301;
  wire [22:0] result_fraction__704;
  wire ne_163380;
  wire ne_163382;
  wire eq_163383;
  wire eq_163384;
  wire eq_163385;
  wire eq_163386;
  wire ne_163389;
  wire ne_163391;
  wire eq_163392;
  wire eq_163393;
  wire eq_163394;
  wire eq_163395;
  wire ne_163404;
  wire ne_163406;
  wire eq_163407;
  wire eq_163408;
  wire eq_163409;
  wire eq_163410;
  wire ne_163419;
  wire ne_163421;
  wire eq_163422;
  wire eq_163423;
  wire eq_163424;
  wire eq_163425;
  wire ne_163434;
  wire ne_163436;
  wire eq_163437;
  wire eq_163438;
  wire eq_163439;
  wire eq_163440;
  wire [8:0] wide_exponent__38;
  wire has_pos_inf__12;
  wire has_neg_inf__12;
  wire [8:0] wide_exponent__80;
  wire has_pos_inf__26;
  wire has_neg_inf__26;
  wire [8:0] wide_exponent__137;
  wire has_pos_inf__45;
  wire has_neg_inf__45;
  wire [8:0] wide_exponent__194;
  wire has_pos_inf__64;
  wire has_neg_inf__64;
  wire [31:0] array_index_163484;
  wire [8:0] wide_exponent__12;
  wire has_pos_inf__4;
  wire has_neg_inf__4;
  wire [8:0] wide_exponent__81;
  wire has_pos_inf__27;
  wire has_neg_inf__27;
  wire [8:0] wide_exponent__138;
  wire has_pos_inf__46;
  wire has_neg_inf__46;
  wire [8:0] wide_exponent__195;
  wire has_pos_inf__65;
  wire has_neg_inf__65;
  wire [7:0] x_bexp__503;
  wire [7:0] high_exp__303;
  wire is_result_nan__25;
  wire is_operand_inf__12;
  wire and_reduce_163539;
  wire is_result_nan__54;
  wire is_operand_inf__26;
  wire and_reduce_163552;
  wire is_result_nan__93;
  wire is_operand_inf__45;
  wire and_reduce_163565;
  wire is_result_nan__132;
  wire is_operand_inf__64;
  wire and_reduce_163578;
  wire is_result_nan__134;
  wire is_result_nan__8;
  wire is_operand_inf__4;
  wire and_reduce_163585;
  wire [2:0] fraction_shift__372;
  wire [2:0] fraction_shift__239;
  wire [7:0] high_exp__102;
  wire is_result_nan__55;
  wire is_operand_inf__27;
  wire and_reduce_163596;
  wire [2:0] fraction_shift__390;
  wire [2:0] fraction_shift__274;
  wire [7:0] high_exp__166;
  wire is_result_nan__94;
  wire is_operand_inf__46;
  wire and_reduce_163607;
  wire [2:0] fraction_shift__408;
  wire [2:0] fraction_shift__309;
  wire [7:0] high_exp__232;
  wire is_result_nan__133;
  wire is_operand_inf__65;
  wire and_reduce_163618;
  wire [2:0] fraction_shift__426;
  wire [2:0] fraction_shift__344;
  wire [7:0] high_exp__302;
  wire [7:0] result_exp__209;
  wire [2:0] fraction_shift__373;
  wire [2:0] fraction_shift__240;
  wire [7:0] high_exp__103;
  wire [2:0] fraction_shift__39;
  wire result_sign__422;
  wire [7:0] result_exponent__13;
  wire [2:0] fraction_shift__391;
  wire [2:0] fraction_shift__275;
  wire [7:0] high_exp__167;
  wire [2:0] fraction_shift__80;
  wire result_sign__517;
  wire [7:0] result_exponent__26;
  wire [2:0] fraction_shift__409;
  wire [2:0] fraction_shift__310;
  wire [7:0] high_exp__233;
  wire [2:0] fraction_shift__137;
  wire result_sign__614;
  wire [7:0] result_exponent__45;
  wire [2:0] fraction_shift__427;
  wire [2:0] fraction_shift__345;
  wire [7:0] high_exp__304;
  wire [2:0] fraction_shift__194;
  wire result_sign__720;
  wire [7:0] result_exponent__64;
  wire result_sign__721;
  wire [2:0] fraction_shift__12;
  wire result_sign__423;
  wire [7:0] result_exponent__4;
  wire [27:0] shrl_163667;
  wire [2:0] fraction_shift__81;
  wire result_sign__518;
  wire [7:0] result_exponent__27;
  wire [27:0] shrl_163674;
  wire [2:0] fraction_shift__138;
  wire result_sign__615;
  wire [7:0] result_exponent__46;
  wire [27:0] shrl_163681;
  wire [2:0] fraction_shift__195;
  wire result_sign__722;
  wire [7:0] result_exponent__65;
  wire [27:0] shrl_163688;
  wire [8:0] concat_163691;
  wire [27:0] shrl_163692;
  wire [22:0] result_fraction__75;
  wire [8:0] sum__13;
  wire [27:0] shrl_163698;
  wire [22:0] result_fraction__160;
  wire [8:0] sum__28;
  wire [27:0] shrl_163704;
  wire [22:0] result_fraction__277;
  wire [8:0] sum__47;
  wire [27:0] shrl_163710;
  wire [22:0] result_fraction__394;
  wire [8:0] sum__66;
  wire [22:0] result_fraction__22;
  wire [8:0] sum__5;
  wire [22:0] result_fraction__76;
  wire [22:0] nan_fraction__89;
  wire [22:0] result_fraction__161;
  wire [8:0] sum__29;
  wire [22:0] result_fraction__162;
  wire [22:0] nan_fraction__115;
  wire [22:0] result_fraction__278;
  wire [8:0] sum__48;
  wire [22:0] result_fraction__279;
  wire [22:0] nan_fraction__143;
  wire [22:0] result_fraction__395;
  wire [8:0] sum__67;
  wire [22:0] result_fraction__396;
  wire [22:0] nan_fraction__172;
  wire [22:0] result_fraction__23;
  wire [22:0] nan_fraction__90;
  wire [22:0] result_fraction__77;
  wire [7:0] prod_bexp__54;
  wire [7:0] x_bexp__726;
  wire [22:0] result_fraction__163;
  wire [22:0] nan_fraction__116;
  wire [22:0] result_fraction__164;
  wire [7:0] prod_bexp__107;
  wire [7:0] x_bexp__727;
  wire [22:0] result_fraction__280;
  wire [22:0] nan_fraction__144;
  wire [22:0] result_fraction__281;
  wire [7:0] prod_bexp__179;
  wire [7:0] x_bexp__728;
  wire [22:0] result_fraction__397;
  wire [22:0] nan_fraction__173;
  wire [22:0] result_fraction__398;
  wire [22:0] result_fraction__476;
  wire [7:0] prod_bexp__251;
  wire [7:0] x_bexp__729;
  wire [22:0] result_fraction__24;
  wire [7:0] prod_bexp__18;
  wire [7:0] x_bexp__730;
  wire fraction_is_zero__12;
  wire [22:0] prod_fraction__39;
  wire [7:0] incremented_sum__84;
  wire [22:0] result_fraction__165;
  wire [7:0] prod_bexp__108;
  wire [7:0] x_bexp__731;
  wire fraction_is_zero__26;
  wire [22:0] prod_fraction__79;
  wire [7:0] incremented_sum__102;
  wire [22:0] result_fraction__282;
  wire [7:0] prod_bexp__180;
  wire [7:0] x_bexp__732;
  wire fraction_is_zero__45;
  wire [22:0] prod_fraction__133;
  wire [7:0] incremented_sum__120;
  wire [22:0] result_fraction__399;
  wire [7:0] prod_bexp__252;
  wire [7:0] x_bexp__733;
  wire fraction_is_zero__64;
  wire [22:0] prod_fraction__187;
  wire [7:0] incremented_sum__138;
  wire fraction_is_zero__4;
  wire [22:0] prod_fraction__13;
  wire [7:0] incremented_sum__85;
  wire [27:0] wide_y__26;
  wire [7:0] x_bexpbs_difference__14;
  wire fraction_is_zero__27;
  wire [22:0] prod_fraction__80;
  wire [7:0] incremented_sum__103;
  wire [27:0] wide_y__55;
  wire [7:0] x_bexpbs_difference__27;
  wire fraction_is_zero__46;
  wire [22:0] prod_fraction__134;
  wire [7:0] incremented_sum__121;
  wire [27:0] wide_y__93;
  wire [7:0] x_bexpbs_difference__45;
  wire fraction_is_zero__65;
  wire [22:0] prod_fraction__188;
  wire [7:0] incremented_sum__139;
  wire [27:0] wide_y__131;
  wire [7:0] x_bexpbs_difference__63;
  wire [27:0] wide_y__9;
  wire [7:0] x_bexpbs_difference__5;
  wire [2:0] concat_163907;
  wire [7:0] x_bexp__110;
  wire [7:0] x_bexp__734;
  wire [27:0] wide_y__27;
  wire [7:0] sub_163913;
  wire [27:0] wide_y__56;
  wire [7:0] x_bexpbs_difference__28;
  wire [2:0] concat_163919;
  wire [7:0] x_bexp__219;
  wire [7:0] x_bexp__735;
  wire [27:0] wide_y__57;
  wire [7:0] sub_163925;
  wire [27:0] wide_y__94;
  wire [7:0] x_bexpbs_difference__46;
  wire [2:0] concat_163931;
  wire [7:0] x_bexp__363;
  wire [7:0] x_bexp__736;
  wire [27:0] wide_y__95;
  wire [7:0] sub_163937;
  wire [27:0] wide_y__132;
  wire [7:0] x_bexpbs_difference__64;
  wire [2:0] concat_163943;
  wire [7:0] x_bexp__507;
  wire [7:0] x_bexp__737;
  wire [27:0] wide_y__133;
  wire [7:0] sub_163949;
  wire [2:0] concat_163950;
  wire [7:0] x_bexp__38;
  wire [7:0] x_bexp__738;
  wire [27:0] wide_y__10;
  wire [7:0] sub_163956;
  wire result_sign__62;
  wire [22:0] x_fraction__110;
  wire [27:0] dropped__13;
  wire [2:0] concat_163964;
  wire [7:0] x_bexp__220;
  wire [7:0] x_bexp__739;
  wire [27:0] wide_y__58;
  wire [7:0] sub_163970;
  wire result_sign__132;
  wire [22:0] x_fraction__219;
  wire [27:0] dropped__28;
  wire [2:0] concat_163978;
  wire [7:0] x_bexp__364;
  wire [7:0] x_bexp__740;
  wire [27:0] wide_y__96;
  wire [7:0] sub_163984;
  wire result_sign__229;
  wire [22:0] x_fraction__363;
  wire [27:0] dropped__47;
  wire [2:0] concat_163992;
  wire [7:0] x_bexp__508;
  wire [7:0] x_bexp__741;
  wire [27:0] wide_y__134;
  wire [7:0] sub_163998;
  wire [7:0] high_exp__488;
  wire result_sign__326;
  wire [22:0] x_fraction__507;
  wire [27:0] dropped__66;
  wire result_sign__18;
  wire [22:0] x_fraction__38;
  wire [27:0] dropped__5;
  wire result_sign__63;
  wire [27:0] wide_x__26;
  wire result_sign__133;
  wire [22:0] x_fraction__220;
  wire [27:0] dropped__29;
  wire result_sign__134;
  wire [27:0] wide_x__55;
  wire result_sign__230;
  wire [22:0] x_fraction__364;
  wire [27:0] dropped__48;
  wire result_sign__231;
  wire [27:0] wide_x__93;
  wire result_sign__327;
  wire [22:0] x_fraction__508;
  wire [27:0] dropped__67;
  wire x_sign__125;
  wire result_sign__328;
  wire [27:0] wide_x__131;
  wire result_sign__19;
  wire [27:0] wide_x__9;
  wire result_sign__64;
  wire [27:0] wide_x__27;
  wire result_sign__135;
  wire [27:0] wide_x__56;
  wire result_sign__136;
  wire [27:0] wide_x__57;
  wire result_sign__232;
  wire [27:0] wide_x__94;
  wire result_sign__233;
  wire [27:0] wide_x__95;
  wire result_sign__329;
  wire [27:0] wide_x__132;
  wire result_sign__334;
  wire result_sign__330;
  wire [27:0] wide_x__133;
  wire result_sign__20;
  wire [27:0] wide_x__10;
  wire x_sign__28;
  wire prod_sign__13;
  wire [27:0] neg_164108;
  wire [27:0] sticky__41;
  wire result_sign__137;
  wire [27:0] wide_x__58;
  wire x_sign__55;
  wire prod_sign__27;
  wire [27:0] neg_164117;
  wire [27:0] sticky__88;
  wire result_sign__234;
  wire [27:0] wide_x__96;
  wire x_sign__91;
  wire prod_sign__45;
  wire [27:0] neg_164126;
  wire [27:0] sticky__147;
  wire result_sign__331;
  wire [27:0] wide_x__134;
  wire x_sign__127;
  wire prod_sign__63;
  wire [27:0] neg_164135;
  wire [27:0] sticky__206;
  wire x_sign__10;
  wire prod_sign__5;
  wire [27:0] neg_164140;
  wire [27:0] sticky__15;
  wire [27:0] xddend_y__13;
  wire x_sign__56;
  wire prod_sign__28;
  wire [27:0] neg_164149;
  wire [27:0] sticky__89;
  wire [27:0] xddend_y__27;
  wire x_sign__92;
  wire prod_sign__46;
  wire [27:0] neg_164158;
  wire [27:0] sticky__148;
  wire [27:0] xddend_y__45;
  wire x_sign__128;
  wire prod_sign__64;
  wire [27:0] neg_164167;
  wire [27:0] sticky__207;
  wire [27:0] xddend_y__63;
  wire [27:0] xddend_y__5;
  wire [24:0] sel_164178;
  wire result_sign__1015;
  wire [27:0] xddend_y__28;
  wire [24:0] sel_164185;
  wire result_sign__1016;
  wire [27:0] xddend_y__46;
  wire [24:0] sel_164192;
  wire result_sign__1017;
  wire [27:0] xddend_y__64;
  wire [24:0] sel_164199;
  wire result_sign__1018;
  wire [24:0] sel_164202;
  wire result_sign__1019;
  wire [24:0] sel_164207;
  wire result_sign__1020;
  wire [24:0] sel_164212;
  wire result_sign__1021;
  wire [24:0] sel_164217;
  wire result_sign__1022;
  wire [25:0] add_164224;
  wire [25:0] add_164227;
  wire [25:0] add_164230;
  wire [25:0] add_164233;
  wire [25:0] add_164234;
  wire [25:0] add_164237;
  wire [25:0] add_164240;
  wire [25:0] add_164243;
  wire [27:0] concat_164248;
  wire [27:0] concat_164251;
  wire [27:0] concat_164254;
  wire [27:0] concat_164257;
  wire [27:0] concat_164258;
  wire [27:0] concat_164261;
  wire [27:0] concat_164264;
  wire [27:0] concat_164267;
  wire [27:0] xbs_fraction__13;
  wire [27:0] xbs_fraction__27;
  wire [27:0] xbs_fraction__45;
  wire [27:0] xbs_fraction__63;
  wire [27:0] xbs_fraction__5;
  wire [27:0] reverse_164283;
  wire [27:0] xbs_fraction__28;
  wire [27:0] reverse_164285;
  wire [27:0] xbs_fraction__46;
  wire [27:0] reverse_164287;
  wire [27:0] xbs_fraction__64;
  wire [27:0] reverse_164289;
  wire [27:0] reverse_164290;
  wire [28:0] one_hot_164291;
  wire [27:0] reverse_164292;
  wire [28:0] one_hot_164293;
  wire [27:0] reverse_164294;
  wire [28:0] one_hot_164295;
  wire [27:0] reverse_164296;
  wire [28:0] one_hot_164297;
  wire [28:0] one_hot_164298;
  wire [4:0] encode_164299;
  wire [28:0] one_hot_164300;
  wire [4:0] encode_164301;
  wire [28:0] one_hot_164302;
  wire [4:0] encode_164303;
  wire [28:0] one_hot_164304;
  wire [4:0] encode_164305;
  wire [4:0] encode_164306;
  wire [4:0] encode_164308;
  wire [4:0] encode_164310;
  wire [4:0] encode_164312;
  wire cancel__14;
  wire carry_bit__13;
  wire [22:0] result_fraction__502;
  wire cancel__28;
  wire carry_bit__28;
  wire [22:0] result_fraction__569;
  wire cancel__47;
  wire carry_bit__47;
  wire [22:0] result_fraction__634;
  wire cancel__66;
  wire carry_bit__66;
  wire [22:0] result_fraction__707;
  wire cancel__5;
  wire carry_bit__5;
  wire [22:0] result_fraction__503;
  wire [27:0] leading_zeroes__13;
  wire cancel__29;
  wire carry_bit__29;
  wire [22:0] result_fraction__570;
  wire [27:0] leading_zeroes__28;
  wire cancel__48;
  wire carry_bit__48;
  wire [22:0] result_fraction__635;
  wire [27:0] leading_zeroes__47;
  wire cancel__67;
  wire carry_bit__67;
  wire [22:0] result_fraction__708;
  wire [27:0] leading_zeroes__66;
  wire [27:0] leading_zeroes__5;
  wire [26:0] carry_fraction__26;
  wire [27:0] add_164379;
  wire [27:0] leading_zeroes__29;
  wire [26:0] carry_fraction__55;
  wire [27:0] add_164392;
  wire [27:0] leading_zeroes__48;
  wire [26:0] carry_fraction__93;
  wire [27:0] add_164405;
  wire [27:0] leading_zeroes__67;
  wire [31:0] array_index_164412;
  wire [26:0] carry_fraction__131;
  wire [27:0] add_164419;
  wire [26:0] carry_fraction__9;
  wire [27:0] add_164426;
  wire [2:0] concat_164427;
  wire [26:0] carry_fraction__27;
  wire [26:0] cancel_fraction__13;
  wire [26:0] carry_fraction__56;
  wire [27:0] add_164436;
  wire [2:0] concat_164437;
  wire [26:0] carry_fraction__57;
  wire [26:0] cancel_fraction__28;
  wire [26:0] carry_fraction__94;
  wire [27:0] add_164446;
  wire [2:0] concat_164447;
  wire [26:0] carry_fraction__95;
  wire [26:0] cancel_fraction__47;
  wire [26:0] carry_fraction__132;
  wire [27:0] add_164456;
  wire [7:0] x_bexp__510;
  wire [2:0] concat_164458;
  wire [26:0] carry_fraction__133;
  wire [26:0] cancel_fraction__66;
  wire [2:0] concat_164461;
  wire [26:0] carry_fraction__10;
  wire [26:0] cancel_fraction__5;
  wire [26:0] shifted_fraction__13;
  wire [2:0] concat_164465;
  wire [26:0] carry_fraction__58;
  wire [26:0] cancel_fraction__29;
  wire result_sign__1023;
  wire [26:0] shifted_fraction__28;
  wire [2:0] concat_164471;
  wire [26:0] carry_fraction__96;
  wire [26:0] cancel_fraction__48;
  wire result_sign__1024;
  wire [26:0] shifted_fraction__47;
  wire [2:0] concat_164477;
  wire [26:0] carry_fraction__134;
  wire [26:0] cancel_fraction__67;
  wire result_sign__1025;
  wire [26:0] shifted_fraction__66;
  wire [26:0] shifted_fraction__5;
  wire result_sign__1026;
  wire [26:0] shifted_fraction__29;
  wire result_sign__1027;
  wire [26:0] shifted_fraction__48;
  wire result_sign__1028;
  wire [26:0] shifted_fraction__67;
  wire result_sign__1029;
  wire result_sign__1030;
  wire [2:0] normal_chunk__13;
  wire [2:0] fraction_shift__241;
  wire [1:0] half_way_chunk__13;
  wire result_sign__1031;
  wire result_sign__1107;
  wire [1:0] add_164512;
  wire [2:0] normal_chunk__28;
  wire [2:0] fraction_shift__276;
  wire [1:0] half_way_chunk__28;
  wire result_sign__1032;
  wire result_sign__1110;
  wire [1:0] add_164523;
  wire [7:0] x_bexp__742;
  wire result_sign__616;
  wire [22:0] x_fraction__505;
  wire [2:0] normal_chunk__47;
  wire [2:0] fraction_shift__311;
  wire [1:0] half_way_chunk__47;
  wire result_sign__1033;
  wire result_sign__1114;
  wire [1:0] add_164537;
  wire [7:0] x_bexp__743;
  wire result_sign__723;
  wire [22:0] x_fraction__510;
  wire [2:0] normal_chunk__66;
  wire [2:0] fraction_shift__346;
  wire [1:0] half_way_chunk__66;
  wire [2:0] normal_chunk__5;
  wire [2:0] fraction_shift__242;
  wire [1:0] half_way_chunk__5;
  wire result_sign__424;
  wire [24:0] add_164557;
  wire [2:0] normal_chunk__29;
  wire [2:0] fraction_shift__277;
  wire [1:0] half_way_chunk__29;
  wire result_sign__519;
  wire [24:0] add_164569;
  wire [2:0] normal_chunk__48;
  wire [2:0] fraction_shift__312;
  wire [1:0] half_way_chunk__48;
  wire ne_164578;
  wire result_sign__618;
  wire [24:0] add_164584;
  wire [2:0] normal_chunk__67;
  wire [2:0] fraction_shift__347;
  wire [1:0] half_way_chunk__67;
  wire ne_164593;
  wire result_sign__725;
  wire [24:0] add_164599;
  wire result_sign__425;
  wire [24:0] add_164603;
  wire do_round_up__27;
  wire result_sign__520;
  wire [24:0] add_164610;
  wire [9:0] exp__124;
  wire do_round_up__58;
  wire result_sign__619;
  wire [24:0] add_164618;
  wire [9:0] exp__206;
  wire [9:0] sign_ext_164620;
  wire [23:0] x_fraction__368;
  wire do_round_up__97;
  wire result_sign__726;
  wire [24:0] add_164629;
  wire [9:0] exp__288;
  wire [9:0] sign_ext_164631;
  wire [23:0] x_fraction__512;
  wire do_round_up__136;
  wire do_round_up__10;
  wire [27:0] rounded_fraction__13;
  wire do_round_up__59;
  wire [9:0] exp__126;
  wire [27:0] rounded_fraction__28;
  wire do_round_up__98;
  wire [9:0] exp__208;
  wire [23:0] x_fraction__370;
  wire result_sign__816;
  wire result_sign__817;
  wire [27:0] rounded_fraction__47;
  wire do_round_up__137;
  wire [9:0] exp__290;
  wire [23:0] x_fraction__514;
  wire result_sign__818;
  wire result_sign__819;
  wire [27:0] rounded_fraction__66;
  wire [27:0] rounded_fraction__5;
  wire result_sign__426;
  wire [7:0] x_bexp__582;
  wire rounding_carry__13;
  wire [27:0] rounded_fraction__29;
  wire result_sign__521;
  wire [7:0] x_bexp__600;
  wire rounding_carry__28;
  wire [27:0] rounded_fraction__48;
  wire [24:0] concat_164676;
  wire [24:0] concat_164677;
  wire result_sign__620;
  wire [7:0] x_bexp__618;
  wire rounding_carry__47;
  wire [27:0] rounded_fraction__67;
  wire [24:0] concat_164683;
  wire [24:0] concat_164684;
  wire result_sign__727;
  wire [7:0] x_bexp__636;
  wire rounding_carry__66;
  wire result_sign__427;
  wire [7:0] x_bexp__583;
  wire rounding_carry__5;
  wire result_sign__522;
  wire [7:0] x_bexp__601;
  wire rounding_carry__29;
  wire [24:0] sel_164696;
  wire result_sign__621;
  wire [7:0] x_bexp__619;
  wire rounding_carry__48;
  wire [24:0] sel_164702;
  wire result_sign__728;
  wire [7:0] x_bexp__637;
  wire rounding_carry__67;
  wire [24:0] sel_164708;
  wire result_sign__428;
  wire [8:0] add_164714;
  wire result_sign__937;
  wire [22:0] fraction__281;
  wire result_sign__523;
  wire [8:0] add_164722;
  wire result_sign__944;
  wire [22:0] fraction__460;
  wire result_sign__622;
  wire [8:0] add_164730;
  wire result_sign__952;
  wire [22:0] fraction__639;
  wire result_sign__729;
  wire [8:0] add_164738;
  wire result_sign__429;
  wire [8:0] add_164742;
  wire result_sign__524;
  wire [8:0] add_164751;
  wire [23:0] fraction__283;
  wire result_sign__623;
  wire [8:0] add_164764;
  wire [23:0] fraction__462;
  wire result_sign__730;
  wire [8:0] add_164777;
  wire [23:0] fraction__641;
  wire [9:0] add_164794;
  wire do_round_up__61;
  wire [23:0] add_164803;
  wire [9:0] add_164804;
  wire do_round_up__100;
  wire [23:0] add_164813;
  wire [9:0] add_164814;
  wire do_round_up__139;
  wire [23:0] add_164823;
  wire [9:0] add_164824;
  wire [9:0] add_164827;
  wire [9:0] wide_exponent__39;
  wire [9:0] add_164832;
  wire [23:0] fraction__285;
  wire [9:0] wide_exponent__82;
  wire [9:0] add_164839;
  wire [23:0] fraction__464;
  wire [9:0] wide_exponent__139;
  wire [9:0] add_164846;
  wire [23:0] fraction__643;
  wire [9:0] wide_exponent__196;
  wire [9:0] wide_exponent__13;
  wire [9:0] wide_exponent__40;
  wire [9:0] wide_exponent__83;
  wire [9:0] add_164859;
  wire [9:0] wide_exponent__84;
  wire [9:0] wide_exponent__140;
  wire [9:0] add_164864;
  wire [9:0] wide_exponent__141;
  wire [9:0] wide_exponent__197;
  wire [9:0] add_164869;
  wire [9:0] wide_exponent__198;
  wire [9:0] wide_exponent__14;
  wire [7:0] high_exp__371;
  wire [22:0] result_fraction__777;
  wire [7:0] high_exp__372;
  wire [22:0] result_fraction__778;
  wire [7:0] high_exp__104;
  wire [22:0] result_fraction__504;
  wire [7:0] high_exp__105;
  wire [22:0] result_fraction__505;
  wire [9:0] wide_exponent__85;
  wire [9:0] exp__130;
  wire [7:0] high_exp__403;
  wire [22:0] result_fraction__810;
  wire [7:0] high_exp__404;
  wire [22:0] result_fraction__811;
  wire [7:0] high_exp__168;
  wire [22:0] result_fraction__571;
  wire [7:0] high_exp__169;
  wire [22:0] result_fraction__572;
  wire [9:0] wide_exponent__142;
  wire [9:0] exp__212;
  wire [7:0] high_exp__435;
  wire [22:0] result_fraction__843;
  wire [7:0] high_exp__436;
  wire [22:0] result_fraction__844;
  wire [7:0] high_exp__234;
  wire [22:0] result_fraction__636;
  wire [7:0] high_exp__235;
  wire [22:0] result_fraction__637;
  wire [9:0] wide_exponent__199;
  wire [9:0] exp__294;
  wire [7:0] high_exp__467;
  wire [22:0] result_fraction__876;
  wire [7:0] high_exp__468;
  wire [22:0] result_fraction__877;
  wire [7:0] high_exp__305;
  wire [22:0] result_fraction__709;
  wire [7:0] high_exp__306;
  wire [22:0] result_fraction__710;
  wire [7:0] high_exp__357;
  wire [22:0] result_fraction__762;
  wire [7:0] high_exp__358;
  wire [22:0] result_fraction__763;
  wire [7:0] high_exp__106;
  wire [22:0] result_fraction__506;
  wire [7:0] high_exp__107;
  wire [22:0] result_fraction__507;
  wire ne_164928;
  wire ne_164930;
  wire eq_164931;
  wire eq_164932;
  wire eq_164933;
  wire eq_164934;
  wire [7:0] high_exp__389;
  wire [22:0] result_fraction__795;
  wire [7:0] high_exp__390;
  wire [22:0] result_fraction__796;
  wire [7:0] high_exp__170;
  wire [22:0] result_fraction__573;
  wire [7:0] high_exp__171;
  wire [22:0] result_fraction__574;
  wire ne_164947;
  wire ne_164949;
  wire eq_164950;
  wire eq_164951;
  wire eq_164952;
  wire eq_164953;
  wire [7:0] high_exp__421;
  wire [22:0] result_fraction__828;
  wire [7:0] high_exp__422;
  wire [22:0] result_fraction__829;
  wire [7:0] high_exp__236;
  wire [22:0] result_fraction__638;
  wire [7:0] high_exp__237;
  wire [22:0] result_fraction__639;
  wire ne_164966;
  wire ne_164968;
  wire eq_164969;
  wire eq_164970;
  wire eq_164971;
  wire eq_164972;
  wire [7:0] high_exp__453;
  wire [22:0] result_fraction__861;
  wire [7:0] high_exp__454;
  wire [22:0] result_fraction__862;
  wire [7:0] high_exp__307;
  wire [22:0] result_fraction__711;
  wire [7:0] high_exp__308;
  wire [22:0] result_fraction__712;
  wire ne_164985;
  wire ne_164987;
  wire eq_164988;
  wire eq_164989;
  wire eq_164990;
  wire eq_164991;
  wire ne_164994;
  wire ne_164996;
  wire eq_164997;
  wire eq_164998;
  wire eq_164999;
  wire eq_165000;
  wire ne_165009;
  wire ne_165011;
  wire eq_165012;
  wire eq_165013;
  wire eq_165014;
  wire eq_165015;
  wire [8:0] result_exp__92;
  wire ne_165026;
  wire ne_165028;
  wire eq_165029;
  wire eq_165030;
  wire eq_165031;
  wire eq_165032;
  wire [8:0] result_exp__152;
  wire ne_165043;
  wire ne_165045;
  wire eq_165046;
  wire eq_165047;
  wire eq_165048;
  wire eq_165049;
  wire [8:0] result_exp__212;
  wire [8:0] wide_exponent__41;
  wire has_pos_inf__13;
  wire has_neg_inf__13;
  wire [8:0] result_exp__94;
  wire [8:0] wide_exponent__86;
  wire has_pos_inf__28;
  wire has_neg_inf__28;
  wire [22:0] result_fraction__706;
  wire [22:0] result_fraction__705;
  wire [8:0] result_exp__154;
  wire [8:0] wide_exponent__143;
  wire has_pos_inf__47;
  wire has_neg_inf__47;
  wire [7:0] high_exp__310;
  wire [22:0] result_fraction__714;
  wire [22:0] result_fraction__713;
  wire [8:0] result_exp__214;
  wire [8:0] wide_exponent__200;
  wire has_pos_inf__66;
  wire has_neg_inf__66;
  wire [8:0] wide_exponent__15;
  wire has_pos_inf__5;
  wire has_neg_inf__5;
  wire [8:0] wide_exponent__87;
  wire has_pos_inf__29;
  wire has_neg_inf__29;
  wire [8:0] wide_exponent__144;
  wire has_pos_inf__48;
  wire has_neg_inf__48;
  wire ne_165126;
  wire [8:0] wide_exponent__201;
  wire has_pos_inf__67;
  wire has_neg_inf__67;
  wire is_result_nan__138;
  wire ne_165140;
  wire is_result_nan__27;
  wire is_operand_inf__13;
  wire and_reduce_165162;
  wire and_reduce_165171;
  wire is_result_nan__58;
  wire is_operand_inf__28;
  wire and_reduce_165177;
  wire is_result_nan__100;
  wire has_inf_arg__69;
  wire and_reduce_165188;
  wire is_result_nan__97;
  wire is_operand_inf__47;
  wire and_reduce_165194;
  wire is_result_nan__139;
  wire has_inf_arg__71;
  wire and_reduce_165205;
  wire is_result_nan__136;
  wire is_operand_inf__66;
  wire and_reduce_165211;
  wire is_result_nan__10;
  wire is_operand_inf__5;
  wire and_reduce_165217;
  wire [2:0] fraction_shift__374;
  wire [2:0] fraction_shift__243;
  wire [7:0] high_exp__108;
  wire is_result_nan__59;
  wire is_operand_inf__29;
  wire and_reduce_165229;
  wire [7:0] high_exp__174;
  wire [2:0] fraction_shift__392;
  wire [2:0] fraction_shift__278;
  wire [7:0] high_exp__172;
  wire [7:0] result_exp__95;
  wire is_result_nan__98;
  wire is_operand_inf__48;
  wire and_reduce_165244;
  wire [7:0] high_exp__240;
  wire [2:0] fraction_shift__410;
  wire [2:0] fraction_shift__313;
  wire [7:0] high_exp__238;
  wire is_result_nan__137;
  wire is_operand_inf__67;
  wire and_reduce_165258;
  wire [7:0] high_exp__312;
  wire [2:0] fraction_shift__428;
  wire [2:0] fraction_shift__348;
  wire [7:0] high_exp__309;
  wire [7:0] result_exp__215;
  wire [2:0] fraction_shift__375;
  wire [2:0] fraction_shift__244;
  wire [7:0] high_exp__109;
  wire [2:0] fraction_shift__42;
  wire result_sign__430;
  wire [7:0] result_exponent__14;
  wire [2:0] fraction_shift__393;
  wire [2:0] fraction_shift__279;
  wire is_subnormal__32;
  wire [7:0] high_exp__173;
  wire [7:0] result_exp__96;
  wire [2:0] fraction_shift__86;
  wire result_sign__525;
  wire [7:0] result_exponent__28;
  wire result_sign__526;
  wire [2:0] fraction_shift__411;
  wire [2:0] fraction_shift__314;
  wire is_subnormal__52;
  wire [7:0] high_exp__239;
  wire [7:0] result_exp__156;
  wire [2:0] fraction_shift__143;
  wire result_sign__624;
  wire [7:0] result_exponent__47;
  wire [2:0] fraction_shift__429;
  wire [2:0] fraction_shift__349;
  wire is_subnormal__72;
  wire [7:0] high_exp__311;
  wire [7:0] result_exp__216;
  wire [2:0] fraction_shift__200;
  wire result_sign__731;
  wire [7:0] result_exponent__66;
  wire result_sign__732;
  wire [2:0] fraction_shift__15;
  wire result_sign__431;
  wire [7:0] result_exponent__5;
  wire [27:0] shrl_165317;
  wire [2:0] fraction_shift__87;
  wire result_sign__527;
  wire [7:0] result_exponent__29;
  wire result_sign__528;
  wire [27:0] shrl_165327;
  wire [2:0] fraction_shift__144;
  wire result_sign__625;
  wire [7:0] result_exponent__48;
  wire result_sign__626;
  wire [27:0] shrl_165338;
  wire [2:0] fraction_shift__201;
  wire result_sign__733;
  wire [7:0] result_exponent__67;
  wire result_sign__734;
  wire [27:0] shrl_165348;
  wire [27:0] shrl_165352;
  wire [22:0] result_fraction__81;
  wire [8:0] sum__14;
  wire [27:0] shrl_165358;
  wire [22:0] result_fraction__172;
  wire [8:0] sum__30;
  wire [27:0] shrl_165366;
  wire [8:0] concat_165370;
  wire [22:0] result_fraction__289;
  wire [8:0] sum__49;
  wire [27:0] shrl_165374;
  wire [22:0] result_fraction__406;
  wire [8:0] sum__68;
  wire [22:0] result_fraction__28;
  wire [8:0] sum__6;
  wire [22:0] result_fraction__82;
  wire [22:0] nan_fraction__91;
  wire [22:0] result_fraction__173;
  wire [22:0] result_fraction__179;
  wire [8:0] sum__31;
  wire [22:0] result_fraction__174;
  wire [22:0] nan_fraction__117;
  wire [22:0] result_fraction__290;
  wire [22:0] result_fraction__296;
  wire [8:0] sum__50;
  wire [22:0] result_fraction__291;
  wire [22:0] nan_fraction__145;
  wire [22:0] result_fraction__407;
  wire [22:0] result_fraction__413;
  wire [8:0] sum__69;
  wire [22:0] result_fraction__408;
  wire [22:0] nan_fraction__174;
  wire [22:0] result_fraction__29;
  wire [22:0] nan_fraction__92;
  wire [22:0] result_fraction__83;
  wire [7:0] prod_bexp__58;
  wire [7:0] x_bexp__744;
  wire [22:0] result_fraction__175;
  wire [22:0] nan_fraction__118;
  wire [22:0] result_fraction__181;
  wire [22:0] nan_fraction__119;
  wire [22:0] result_fraction__176;
  wire [22:0] result_fraction__477;
  wire [7:0] prod_bexp__115;
  wire [7:0] x_bexp__745;
  wire [22:0] result_fraction__292;
  wire [22:0] nan_fraction__146;
  wire [22:0] result_fraction__298;
  wire [22:0] nan_fraction__147;
  wire [22:0] result_fraction__293;
  wire [7:0] prod_bexp__187;
  wire [7:0] x_bexp__746;
  wire [22:0] result_fraction__409;
  wire [22:0] nan_fraction__175;
  wire [22:0] result_fraction__415;
  wire [22:0] nan_fraction__176;
  wire [22:0] result_fraction__410;
  wire [22:0] result_fraction__478;
  wire [7:0] prod_bexp__259;
  wire [7:0] x_bexp__747;
  wire [22:0] result_fraction__30;
  wire [7:0] prod_bexp__22;
  wire [7:0] x_bexp__748;
  wire fraction_is_zero__13;
  wire [22:0] prod_fraction__42;
  wire [7:0] incremented_sum__86;
  wire [22:0] result_fraction__177;
  wire [22:0] result_fraction__183;
  wire [7:0] prod_bexp__116;
  wire [7:0] x_bexp__749;
  wire fraction_is_zero__28;
  wire [22:0] prod_fraction__85;
  wire [7:0] incremented_sum__104;
  wire [22:0] result_fraction__294;
  wire [22:0] result_fraction__300;
  wire [7:0] prod_bexp__188;
  wire [7:0] x_bexp__750;
  wire fraction_is_zero__47;
  wire [22:0] prod_fraction__139;
  wire [7:0] incremented_sum__122;
  wire [22:0] result_fraction__411;
  wire [22:0] result_fraction__417;
  wire [7:0] prod_bexp__260;
  wire [7:0] x_bexp__751;
  wire fraction_is_zero__66;
  wire [22:0] prod_fraction__193;
  wire [7:0] incremented_sum__140;
  wire fraction_is_zero__5;
  wire [22:0] prod_fraction__16;
  wire [7:0] incremented_sum__87;
  wire [27:0] wide_y__28;
  wire [7:0] x_bexpbs_difference__15;
  wire fraction_is_zero__29;
  wire [22:0] prod_fraction__86;
  wire [7:0] incremented_sum__105;
  wire [27:0] wide_y__59;
  wire [7:0] x_bexpbs_difference__29;
  wire fraction_is_zero__48;
  wire [22:0] prod_fraction__140;
  wire [7:0] incremented_sum__123;
  wire [27:0] wide_y__97;
  wire [7:0] x_bexpbs_difference__47;
  wire fraction_is_zero__67;
  wire [22:0] prod_fraction__194;
  wire [7:0] incremented_sum__141;
  wire [27:0] wide_y__135;
  wire [7:0] x_bexpbs_difference__65;
  wire [27:0] wide_y__11;
  wire [7:0] x_bexpbs_difference__6;
  wire [2:0] concat_165590;
  wire [7:0] x_bexp__118;
  wire [7:0] x_bexp__752;
  wire [27:0] wide_y__29;
  wire [7:0] sub_165596;
  wire [27:0] wide_y__60;
  wire [7:0] x_bexpbs_difference__30;
  wire [2:0] concat_165602;
  wire [7:0] x_bexp__235;
  wire [7:0] x_bexp__753;
  wire [27:0] wide_y__61;
  wire [7:0] sub_165608;
  wire [27:0] wide_y__98;
  wire [7:0] x_bexpbs_difference__48;
  wire [2:0] concat_165614;
  wire [7:0] x_bexp__379;
  wire [7:0] x_bexp__754;
  wire [27:0] wide_y__99;
  wire [7:0] sub_165620;
  wire [27:0] wide_y__136;
  wire [7:0] x_bexpbs_difference__66;
  wire [2:0] concat_165626;
  wire [7:0] x_bexp__523;
  wire [7:0] x_bexp__755;
  wire [27:0] wide_y__137;
  wire [7:0] sub_165632;
  wire [2:0] concat_165633;
  wire [7:0] x_bexp__46;
  wire [7:0] x_bexp__756;
  wire [27:0] wide_y__12;
  wire [7:0] sub_165639;
  wire result_sign__67;
  wire [22:0] x_fraction__118;
  wire [27:0] dropped__14;
  wire [2:0] concat_165647;
  wire [7:0] x_bexp__236;
  wire [7:0] x_bexp__757;
  wire [27:0] wide_y__62;
  wire [7:0] sub_165653;
  wire [7:0] high_exp__482;
  wire result_sign__142;
  wire [22:0] x_fraction__235;
  wire [27:0] dropped__30;
  wire [2:0] concat_165662;
  wire [7:0] x_bexp__380;
  wire [7:0] x_bexp__758;
  wire [27:0] wide_y__100;
  wire [7:0] sub_165668;
  wire result_sign__239;
  wire [22:0] x_fraction__379;
  wire [27:0] dropped__49;
  wire [2:0] concat_165676;
  wire [7:0] x_bexp__524;
  wire [7:0] x_bexp__759;
  wire [27:0] wide_y__138;
  wire [7:0] sub_165682;
  wire [7:0] high_exp__489;
  wire result_sign__336;
  wire [22:0] x_fraction__523;
  wire [27:0] dropped__68;
  wire result_sign__23;
  wire [22:0] x_fraction__46;
  wire [27:0] dropped__6;
  wire result_sign__68;
  wire [27:0] wide_x__28;
  wire result_sign__143;
  wire [22:0] x_fraction__236;
  wire [27:0] dropped__31;
  wire result_sign__144;
  wire [27:0] wide_x__59;
  wire result_sign__240;
  wire [22:0] x_fraction__380;
  wire [27:0] dropped__50;
  wire result_sign__241;
  wire [27:0] wide_x__97;
  wire result_sign__337;
  wire [22:0] x_fraction__524;
  wire [27:0] dropped__69;
  wire x_sign__129;
  wire result_sign__338;
  wire [27:0] wide_x__135;
  wire result_sign__24;
  wire [27:0] wide_x__11;
  wire result_sign__69;
  wire [27:0] wide_x__29;
  wire result_sign__145;
  wire [27:0] wide_x__60;
  wire result_sign__150;
  wire result_sign__146;
  wire [27:0] wide_x__61;
  wire result_sign__242;
  wire [27:0] wide_x__98;
  wire result_sign__243;
  wire [27:0] wide_x__99;
  wire result_sign__339;
  wire [27:0] wide_x__136;
  wire result_sign__344;
  wire result_sign__340;
  wire [27:0] wide_x__137;
  wire result_sign__25;
  wire [27:0] wide_x__12;
  wire x_sign__30;
  wire prod_sign__14;
  wire [27:0] neg_165796;
  wire [27:0] sticky__44;
  wire result_sign__147;
  wire [27:0] wide_x__62;
  wire x_sign__59;
  wire prod_sign__29;
  wire [27:0] neg_165805;
  wire [27:0] sticky__94;
  wire result_sign__248;
  wire result_sign__244;
  wire [27:0] wide_x__100;
  wire x_sign__95;
  wire prod_sign__47;
  wire [27:0] neg_165815;
  wire [27:0] sticky__153;
  wire result_sign__345;
  wire result_sign__341;
  wire [27:0] wide_x__138;
  wire x_sign__131;
  wire prod_sign__65;
  wire [27:0] neg_165825;
  wire [27:0] sticky__212;
  wire x_sign__12;
  wire prod_sign__6;
  wire [27:0] neg_165830;
  wire [27:0] sticky__18;
  wire [27:0] xddend_y__14;
  wire x_sign__60;
  wire prod_sign__30;
  wire [27:0] neg_165839;
  wire [27:0] sticky__95;
  wire [27:0] xddend_y__29;
  wire x_sign__96;
  wire prod_sign__48;
  wire [27:0] neg_165848;
  wire [27:0] sticky__154;
  wire [27:0] xddend_y__47;
  wire x_sign__132;
  wire prod_sign__66;
  wire [27:0] neg_165857;
  wire [27:0] sticky__213;
  wire [27:0] xddend_y__65;
  wire [27:0] xddend_y__6;
  wire [24:0] sel_165868;
  wire result_sign__1034;
  wire [27:0] xddend_y__30;
  wire [24:0] sel_165875;
  wire result_sign__1035;
  wire [27:0] xddend_y__48;
  wire [24:0] sel_165882;
  wire result_sign__1036;
  wire [27:0] xddend_y__66;
  wire [24:0] sel_165889;
  wire result_sign__1037;
  wire [24:0] sel_165892;
  wire result_sign__1038;
  wire [24:0] sel_165897;
  wire result_sign__1039;
  wire [24:0] sel_165902;
  wire result_sign__1040;
  wire [24:0] sel_165907;
  wire result_sign__1041;
  wire [25:0] add_165914;
  wire [25:0] add_165917;
  wire [25:0] add_165920;
  wire [25:0] add_165923;
  wire [25:0] add_165924;
  wire [25:0] add_165927;
  wire [25:0] add_165930;
  wire [25:0] add_165933;
  wire [27:0] concat_165938;
  wire [27:0] concat_165941;
  wire [27:0] concat_165944;
  wire [27:0] concat_165947;
  wire [27:0] concat_165948;
  wire [27:0] concat_165951;
  wire [27:0] concat_165954;
  wire [27:0] concat_165957;
  wire [27:0] xbs_fraction__14;
  wire [27:0] xbs_fraction__29;
  wire [27:0] xbs_fraction__47;
  wire [27:0] xbs_fraction__65;
  wire [27:0] xbs_fraction__6;
  wire [27:0] reverse_165973;
  wire [27:0] xbs_fraction__30;
  wire [27:0] reverse_165975;
  wire [27:0] xbs_fraction__48;
  wire [27:0] reverse_165977;
  wire [27:0] xbs_fraction__66;
  wire [27:0] reverse_165979;
  wire [27:0] reverse_165980;
  wire [28:0] one_hot_165981;
  wire [27:0] reverse_165982;
  wire [28:0] one_hot_165983;
  wire [27:0] reverse_165984;
  wire [28:0] one_hot_165985;
  wire [27:0] reverse_165986;
  wire [28:0] one_hot_165987;
  wire [28:0] one_hot_165988;
  wire [4:0] encode_165989;
  wire [28:0] one_hot_165990;
  wire [4:0] encode_165991;
  wire [28:0] one_hot_165992;
  wire [4:0] encode_165993;
  wire [28:0] one_hot_165994;
  wire [4:0] encode_165995;
  wire [4:0] encode_165996;
  wire [4:0] encode_165998;
  wire [4:0] encode_166000;
  wire [4:0] encode_166002;
  wire cancel__15;
  wire carry_bit__14;
  wire [22:0] result_fraction__508;
  wire cancel__30;
  wire carry_bit__30;
  wire [22:0] result_fraction__575;
  wire cancel__49;
  wire carry_bit__49;
  wire [22:0] result_fraction__640;
  wire cancel__68;
  wire carry_bit__68;
  wire [22:0] result_fraction__715;
  wire cancel__6;
  wire carry_bit__6;
  wire [22:0] result_fraction__509;
  wire [27:0] leading_zeroes__14;
  wire cancel__31;
  wire carry_bit__31;
  wire [22:0] result_fraction__576;
  wire [27:0] leading_zeroes__30;
  wire cancel__50;
  wire carry_bit__50;
  wire [22:0] result_fraction__641;
  wire [27:0] leading_zeroes__49;
  wire cancel__69;
  wire carry_bit__69;
  wire [22:0] result_fraction__716;
  wire [27:0] leading_zeroes__68;
  wire [27:0] leading_zeroes__6;
  wire [26:0] carry_fraction__28;
  wire [27:0] add_166070;
  wire [27:0] leading_zeroes__31;
  wire [26:0] carry_fraction__59;
  wire [27:0] add_166083;
  wire [27:0] leading_zeroes__50;
  wire [26:0] carry_fraction__97;
  wire [27:0] add_166096;
  wire [31:0] array_index_166097;
  wire [27:0] leading_zeroes__69;
  wire [26:0] carry_fraction__135;
  wire [27:0] add_166110;
  wire [31:0] array_index_166111;
  wire [26:0] carry_fraction__11;
  wire [27:0] add_166118;
  wire [2:0] concat_166119;
  wire [26:0] carry_fraction__29;
  wire [26:0] cancel_fraction__14;
  wire result_sign__599;
  wire [26:0] carry_fraction__60;
  wire [27:0] add_166129;
  wire [2:0] concat_166130;
  wire [26:0] carry_fraction__61;
  wire [26:0] cancel_fraction__30;
  wire result_sign__705;
  wire [26:0] carry_fraction__98;
  wire [27:0] add_166140;
  wire [2:0] concat_166141;
  wire [26:0] carry_fraction__99;
  wire [26:0] cancel_fraction__49;
  wire result_sign__630;
  wire [7:0] x_bexp__381;
  wire [26:0] carry_fraction__136;
  wire [27:0] add_166152;
  wire [2:0] concat_166153;
  wire [26:0] carry_fraction__137;
  wire [26:0] cancel_fraction__68;
  wire result_sign__738;
  wire [7:0] x_bexp__525;
  wire [2:0] concat_166158;
  wire [26:0] carry_fraction__12;
  wire [26:0] cancel_fraction__6;
  wire [26:0] shifted_fraction__14;
  wire [2:0] concat_166164;
  wire [26:0] carry_fraction__62;
  wire [26:0] cancel_fraction__31;
  wire [26:0] shifted_fraction__30;
  wire [2:0] concat_166170;
  wire [26:0] carry_fraction__100;
  wire [26:0] cancel_fraction__50;
  wire [26:0] shifted_fraction__49;
  wire [2:0] concat_166176;
  wire [26:0] carry_fraction__138;
  wire [26:0] cancel_fraction__69;
  wire [26:0] shifted_fraction__68;
  wire [26:0] shifted_fraction__6;
  wire result_sign__1042;
  wire result_sign__435;
  wire [8:0] add_166186;
  wire [26:0] shifted_fraction__31;
  wire result_sign__1043;
  wire result_sign__532;
  wire [8:0] add_166191;
  wire [26:0] shifted_fraction__50;
  wire result_sign__1044;
  wire result_sign__632;
  wire [8:0] add_166196;
  wire [7:0] x_bexp__760;
  wire result_sign__628;
  wire [22:0] x_fraction__381;
  wire [26:0] shifted_fraction__69;
  wire result_sign__1045;
  wire result_sign__740;
  wire [8:0] add_166204;
  wire [7:0] x_bexp__761;
  wire result_sign__736;
  wire [22:0] x_fraction__525;
  wire result_sign__1046;
  wire [2:0] normal_chunk__14;
  wire [2:0] fraction_shift__245;
  wire [1:0] half_way_chunk__14;
  wire result_sign__1047;
  wire [2:0] normal_chunk__30;
  wire [2:0] fraction_shift__280;
  wire [1:0] half_way_chunk__30;
  wire result_sign__1048;
  wire [2:0] normal_chunk__49;
  wire [2:0] fraction_shift__315;
  wire [1:0] half_way_chunk__49;
  wire ne_166238;
  wire result_sign__1049;
  wire [2:0] normal_chunk__68;
  wire [2:0] fraction_shift__350;
  wire [1:0] half_way_chunk__68;
  wire ne_166251;
  wire [2:0] normal_chunk__6;
  wire [2:0] fraction_shift__246;
  wire [1:0] half_way_chunk__6;
  wire result_sign__432;
  wire [24:0] add_166263;
  wire [9:0] exp__60;
  wire [2:0] normal_chunk__31;
  wire [2:0] fraction_shift__281;
  wire [1:0] half_way_chunk__31;
  wire result_sign__529;
  wire [24:0] add_166274;
  wire [9:0] exp__131;
  wire [2:0] normal_chunk__50;
  wire [2:0] fraction_shift__316;
  wire [1:0] half_way_chunk__50;
  wire result_sign__627;
  wire [24:0] add_166285;
  wire [9:0] exp__213;
  wire [23:0] x_fraction__383;
  wire [2:0] normal_chunk__69;
  wire [2:0] fraction_shift__351;
  wire [1:0] half_way_chunk__69;
  wire result_sign__735;
  wire [24:0] add_166299;
  wire [9:0] exp__295;
  wire [9:0] sign_ext_166301;
  wire [23:0] x_fraction__527;
  wire result_sign__433;
  wire [24:0] add_166307;
  wire do_round_up__29;
  wire [9:0] exp__61;
  wire result_sign__530;
  wire [24:0] add_166316;
  wire do_round_up__62;
  wire [9:0] exp__133;
  wire result_sign__629;
  wire [24:0] add_166325;
  wire do_round_up__101;
  wire [9:0] exp__215;
  wire [23:0] x_fraction__385;
  wire result_sign__820;
  wire result_sign__821;
  wire result_sign__737;
  wire [24:0] add_166337;
  wire do_round_up__140;
  wire [9:0] exp__297;
  wire [23:0] x_fraction__529;
  wire result_sign__822;
  wire result_sign__823;
  wire do_round_up__12;
  wire [27:0] rounded_fraction__14;
  wire do_round_up__63;
  wire [27:0] rounded_fraction__30;
  wire do_round_up__102;
  wire [27:0] rounded_fraction__49;
  wire do_round_up__141;
  wire [27:0] rounded_fraction__68;
  wire [24:0] concat_166368;
  wire [24:0] concat_166369;
  wire [27:0] rounded_fraction__6;
  wire result_sign__434;
  wire [7:0] x_bexp__584;
  wire rounding_carry__14;
  wire [24:0] sel_166374;
  wire [27:0] rounded_fraction__31;
  wire result_sign__531;
  wire [7:0] x_bexp__602;
  wire rounding_carry__30;
  wire [24:0] sel_166379;
  wire [27:0] rounded_fraction__50;
  wire result_sign__631;
  wire [7:0] x_bexp__620;
  wire rounding_carry__49;
  wire [24:0] sel_166384;
  wire [27:0] rounded_fraction__69;
  wire result_sign__739;
  wire [7:0] x_bexp__638;
  wire rounding_carry__68;
  wire [24:0] sel_166389;
  wire result_sign__436;
  wire [7:0] x_bexp__585;
  wire rounding_carry__6;
  wire result_sign__932;
  wire [22:0] fraction__140;
  wire result_sign__533;
  wire [7:0] x_bexp__603;
  wire rounding_carry__31;
  wire result_sign__938;
  wire [22:0] fraction__298;
  wire result_sign__633;
  wire [7:0] x_bexp__621;
  wire rounding_carry__50;
  wire result_sign__945;
  wire [22:0] fraction__477;
  wire result_sign__741;
  wire [7:0] x_bexp__639;
  wire rounding_carry__69;
  wire result_sign__953;
  wire [22:0] fraction__656;
  wire result_sign__437;
  wire [8:0] add_166421;
  wire [23:0] fraction__141;
  wire result_sign__534;
  wire [8:0] add_166431;
  wire [23:0] fraction__300;
  wire result_sign__634;
  wire [8:0] add_166441;
  wire [23:0] fraction__479;
  wire result_sign__742;
  wire [8:0] add_166451;
  wire [23:0] fraction__658;
  wire result_sign__438;
  wire [8:0] add_166459;
  wire do_round_up__30;
  wire [23:0] add_166468;
  wire result_sign__535;
  wire [8:0] add_166470;
  wire do_round_up__64;
  wire [23:0] add_166479;
  wire result_sign__635;
  wire [8:0] add_166481;
  wire do_round_up__103;
  wire [23:0] add_166490;
  wire result_sign__743;
  wire [8:0] add_166492;
  wire do_round_up__142;
  wire [23:0] add_166501;
  wire [9:0] add_166507;
  wire [23:0] fraction__142;
  wire [9:0] add_166517;
  wire [23:0] fraction__302;
  wire [9:0] add_166527;
  wire [23:0] fraction__481;
  wire [9:0] add_166537;
  wire [23:0] fraction__660;
  wire [9:0] add_166542;
  wire [9:0] wide_exponent__42;
  wire [9:0] add_166548;
  wire [9:0] add_166549;
  wire [9:0] wide_exponent__88;
  wire [9:0] add_166555;
  wire [9:0] add_166556;
  wire [9:0] wide_exponent__145;
  wire [9:0] add_166562;
  wire [9:0] add_166563;
  wire [9:0] wide_exponent__202;
  wire [9:0] add_166569;
  wire [9:0] wide_exponent__16;
  wire [9:0] wide_exponent__43;
  wire [9:0] exp__63;
  wire [9:0] wide_exponent__89;
  wire [9:0] wide_exponent__90;
  wire [9:0] exp__137;
  wire [9:0] wide_exponent__146;
  wire [9:0] wide_exponent__147;
  wire [9:0] exp__219;
  wire [9:0] wide_exponent__203;
  wire [9:0] wide_exponent__204;
  wire [9:0] exp__301;
  wire [9:0] wide_exponent__17;
  wire [7:0] high_exp__373;
  wire [22:0] result_fraction__779;
  wire [7:0] high_exp__374;
  wire [22:0] result_fraction__780;
  wire [7:0] high_exp__110;
  wire [22:0] result_fraction__510;
  wire [7:0] high_exp__111;
  wire [22:0] result_fraction__511;
  wire [9:0] wide_exponent__91;
  wire [7:0] high_exp__405;
  wire [22:0] result_fraction__812;
  wire [7:0] high_exp__406;
  wire [22:0] result_fraction__813;
  wire [7:0] high_exp__175;
  wire [22:0] result_fraction__577;
  wire [7:0] high_exp__176;
  wire [22:0] result_fraction__578;
  wire [9:0] wide_exponent__148;
  wire [7:0] high_exp__437;
  wire [22:0] result_fraction__845;
  wire [7:0] high_exp__438;
  wire [22:0] result_fraction__846;
  wire [7:0] high_exp__241;
  wire [22:0] result_fraction__642;
  wire [7:0] high_exp__242;
  wire [22:0] result_fraction__643;
  wire [9:0] wide_exponent__205;
  wire [7:0] high_exp__469;
  wire [22:0] result_fraction__878;
  wire [7:0] high_exp__470;
  wire [22:0] result_fraction__879;
  wire [7:0] high_exp__313;
  wire [22:0] result_fraction__717;
  wire [7:0] high_exp__314;
  wire [22:0] result_fraction__718;
  wire [7:0] high_exp__359;
  wire [22:0] result_fraction__764;
  wire [7:0] high_exp__360;
  wire [22:0] result_fraction__765;
  wire [7:0] high_exp__112;
  wire [22:0] result_fraction__512;
  wire [7:0] high_exp__113;
  wire [22:0] result_fraction__513;
  wire ne_166645;
  wire ne_166647;
  wire eq_166648;
  wire eq_166649;
  wire eq_166650;
  wire eq_166651;
  wire [8:0] result_exp__45;
  wire [7:0] high_exp__391;
  wire [22:0] result_fraction__797;
  wire [7:0] high_exp__392;
  wire [22:0] result_fraction__798;
  wire [7:0] high_exp__177;
  wire [22:0] result_fraction__579;
  wire [7:0] high_exp__178;
  wire [22:0] result_fraction__580;
  wire ne_166665;
  wire ne_166667;
  wire eq_166668;
  wire eq_166669;
  wire eq_166670;
  wire eq_166671;
  wire [8:0] result_exp__97;
  wire [7:0] high_exp__423;
  wire [22:0] result_fraction__830;
  wire [7:0] high_exp__424;
  wire [22:0] result_fraction__831;
  wire [7:0] high_exp__243;
  wire [22:0] result_fraction__644;
  wire [7:0] high_exp__244;
  wire [22:0] result_fraction__645;
  wire ne_166685;
  wire ne_166687;
  wire eq_166688;
  wire eq_166689;
  wire eq_166690;
  wire eq_166691;
  wire [8:0] result_exp__157;
  wire [7:0] high_exp__455;
  wire [22:0] result_fraction__863;
  wire [7:0] high_exp__456;
  wire [22:0] result_fraction__864;
  wire [7:0] high_exp__315;
  wire [22:0] result_fraction__719;
  wire [7:0] high_exp__316;
  wire [22:0] result_fraction__720;
  wire ne_166705;
  wire ne_166707;
  wire eq_166708;
  wire eq_166709;
  wire eq_166710;
  wire eq_166711;
  wire [8:0] result_exp__217;
  wire ne_166716;
  wire ne_166718;
  wire eq_166719;
  wire eq_166720;
  wire eq_166721;
  wire eq_166722;
  wire [8:0] result_exp__46;
  wire ne_166732;
  wire ne_166734;
  wire eq_166735;
  wire eq_166736;
  wire eq_166737;
  wire eq_166738;
  wire [8:0] result_exp__99;
  wire ne_166748;
  wire ne_166750;
  wire eq_166751;
  wire eq_166752;
  wire eq_166753;
  wire eq_166754;
  wire [7:0] high_exp__247;
  wire [22:0] result_fraction__647;
  wire [22:0] result_fraction__646;
  wire [8:0] result_exp__159;
  wire ne_166767;
  wire ne_166769;
  wire eq_166770;
  wire eq_166771;
  wire eq_166772;
  wire eq_166773;
  wire [7:0] high_exp__319;
  wire [22:0] result_fraction__722;
  wire [22:0] result_fraction__721;
  wire [8:0] result_exp__219;
  wire [8:0] wide_exponent__44;
  wire has_pos_inf__14;
  wire has_neg_inf__14;
  wire [8:0] wide_exponent__92;
  wire has_pos_inf__30;
  wire has_neg_inf__30;
  wire [8:0] wide_exponent__149;
  wire has_pos_inf__49;
  wire has_neg_inf__49;
  wire eq_166813;
  wire ne_166814;
  wire [8:0] wide_exponent__206;
  wire has_pos_inf__68;
  wire has_neg_inf__68;
  wire is_result_nan__108;
  wire ne_166827;
  wire [8:0] wide_exponent__18;
  wire has_pos_inf__6;
  wire has_neg_inf__6;
  wire and_reduce_166841;
  wire [8:0] wide_exponent__93;
  wire has_pos_inf__31;
  wire has_neg_inf__31;
  wire and_reduce_166853;
  wire [8:0] wide_exponent__150;
  wire has_pos_inf__50;
  wire has_neg_inf__50;
  wire is_result_nan__103;
  wire has_inf_arg__53;
  wire and_reduce_166867;
  wire [8:0] wide_exponent__207;
  wire has_pos_inf__69;
  wire has_neg_inf__69;
  wire is_result_nan__142;
  wire has_inf_arg__73;
  wire and_reduce_166881;
  wire is_result_nan__29;
  wire is_operand_inf__14;
  wire and_reduce_166895;
  wire [7:0] high_exp__116;
  wire is_result_nan__62;
  wire is_operand_inf__30;
  wire and_reduce_166911;
  wire [7:0] high_exp__181;
  wire is_result_nan__101;
  wire is_operand_inf__49;
  wire and_reduce_166927;
  wire [7:0] high_exp__248;
  wire is_result_nan__140;
  wire is_operand_inf__68;
  wire and_reduce_166943;
  wire [7:0] high_exp__320;
  wire is_result_nan__12;
  wire is_operand_inf__6;
  wire and_reduce_166951;
  wire [2:0] fraction_shift__376;
  wire [2:0] fraction_shift__247;
  wire is_subnormal__15;
  wire [7:0] high_exp__114;
  wire [7:0] result_exp__47;
  wire is_result_nan__63;
  wire is_operand_inf__31;
  wire and_reduce_166964;
  wire [2:0] fraction_shift__394;
  wire [2:0] fraction_shift__282;
  wire is_subnormal__33;
  wire [7:0] high_exp__179;
  wire [7:0] result_exp__101;
  wire is_result_nan__102;
  wire is_operand_inf__50;
  wire and_reduce_166977;
  wire [2:0] fraction_shift__412;
  wire [2:0] fraction_shift__317;
  wire is_subnormal__53;
  wire [7:0] high_exp__245;
  wire [7:0] result_exp__161;
  wire is_result_nan__141;
  wire is_operand_inf__69;
  wire and_reduce_166990;
  wire [2:0] fraction_shift__430;
  wire [2:0] fraction_shift__352;
  wire is_subnormal__73;
  wire [7:0] high_exp__317;
  wire [7:0] result_exp__221;
  wire [2:0] fraction_shift__377;
  wire [2:0] fraction_shift__248;
  wire [7:0] high_exp__115;
  wire [2:0] fraction_shift__45;
  wire result_sign__439;
  wire [7:0] result_exponent__15;
  wire result_sign__440;
  wire [2:0] fraction_shift__395;
  wire [2:0] fraction_shift__283;
  wire [7:0] high_exp__180;
  wire [2:0] fraction_shift__92;
  wire result_sign__536;
  wire [7:0] result_exponent__30;
  wire result_sign__537;
  wire [2:0] fraction_shift__413;
  wire [2:0] fraction_shift__318;
  wire [7:0] high_exp__246;
  wire [2:0] fraction_shift__149;
  wire result_sign__636;
  wire [7:0] result_exponent__49;
  wire result_sign__637;
  wire [2:0] fraction_shift__431;
  wire [2:0] fraction_shift__353;
  wire [7:0] high_exp__318;
  wire [2:0] fraction_shift__206;
  wire result_sign__744;
  wire [7:0] result_exponent__68;
  wire result_sign__745;
  wire [2:0] fraction_shift__18;
  wire result_sign__441;
  wire [7:0] result_exponent__6;
  wire [27:0] shrl_167050;
  wire [8:0] concat_167054;
  wire [2:0] fraction_shift__93;
  wire result_sign__538;
  wire [7:0] result_exponent__31;
  wire [27:0] shrl_167059;
  wire [8:0] concat_167063;
  wire [2:0] fraction_shift__150;
  wire result_sign__638;
  wire [7:0] result_exponent__50;
  wire [27:0] shrl_167068;
  wire [8:0] concat_167072;
  wire [2:0] fraction_shift__207;
  wire result_sign__746;
  wire [7:0] result_exponent__69;
  wire [27:0] shrl_167077;
  wire [8:0] concat_167081;
  wire [27:0] shrl_167082;
  wire [22:0] result_fraction__87;
  wire [22:0] result_fraction__90;
  wire [8:0] sum__15;
  wire [27:0] shrl_167090;
  wire [22:0] result_fraction__184;
  wire [22:0] result_fraction__190;
  wire [8:0] sum__32;
  wire [27:0] shrl_167098;
  wire [22:0] result_fraction__301;
  wire [22:0] result_fraction__307;
  wire [8:0] sum__51;
  wire [27:0] shrl_167106;
  wire [22:0] result_fraction__418;
  wire [22:0] result_fraction__424;
  wire [8:0] sum__70;
  wire [22:0] result_fraction__34;
  wire [8:0] sum__7;
  wire [22:0] result_fraction__88;
  wire [22:0] nan_fraction__93;
  wire [22:0] result_fraction__91;
  wire [22:0] nan_fraction__95;
  wire [22:0] result_fraction__185;
  wire [8:0] sum__33;
  wire [22:0] result_fraction__186;
  wire [22:0] nan_fraction__120;
  wire [22:0] result_fraction__192;
  wire [22:0] nan_fraction__122;
  wire [22:0] result_fraction__302;
  wire [8:0] sum__52;
  wire [22:0] result_fraction__303;
  wire [22:0] nan_fraction__148;
  wire [22:0] result_fraction__309;
  wire [22:0] nan_fraction__150;
  wire [22:0] result_fraction__419;
  wire [8:0] sum__71;
  wire [22:0] result_fraction__420;
  wire [22:0] nan_fraction__177;
  wire [22:0] result_fraction__426;
  wire [22:0] nan_fraction__179;
  wire [22:0] result_fraction__35;
  wire [22:0] nan_fraction__94;
  wire [22:0] result_fraction__89;
  wire [22:0] result_fraction__92;
  wire [7:0] prod_bexp__62;
  wire [7:0] x_bexp__762;
  wire [22:0] result_fraction__187;
  wire [22:0] nan_fraction__121;
  wire [22:0] result_fraction__188;
  wire [22:0] result_fraction__194;
  wire [7:0] prod_bexp__123;
  wire [7:0] x_bexp__763;
  wire [22:0] result_fraction__304;
  wire [22:0] nan_fraction__149;
  wire [22:0] result_fraction__305;
  wire [22:0] result_fraction__311;
  wire [7:0] prod_bexp__195;
  wire [7:0] x_bexp__764;
  wire [22:0] result_fraction__421;
  wire [22:0] nan_fraction__178;
  wire [22:0] result_fraction__422;
  wire [22:0] result_fraction__428;
  wire [7:0] prod_bexp__267;
  wire [7:0] x_bexp__765;
  wire [22:0] result_fraction__36;
  wire [7:0] prod_bexp__26;
  wire [7:0] x_bexp__766;
  wire fraction_is_zero__14;
  wire [22:0] prod_fraction__45;
  wire [7:0] incremented_sum__88;
  wire [22:0] result_fraction__189;
  wire [7:0] prod_bexp__124;
  wire [7:0] x_bexp__767;
  wire fraction_is_zero__30;
  wire [22:0] prod_fraction__91;
  wire [7:0] incremented_sum__106;
  wire [22:0] result_fraction__306;
  wire [7:0] prod_bexp__196;
  wire [7:0] x_bexp__768;
  wire fraction_is_zero__49;
  wire [22:0] prod_fraction__145;
  wire [7:0] incremented_sum__124;
  wire [22:0] result_fraction__423;
  wire [7:0] prod_bexp__268;
  wire [7:0] x_bexp__769;
  wire fraction_is_zero__68;
  wire [22:0] prod_fraction__199;
  wire [7:0] incremented_sum__142;
  wire fraction_is_zero__6;
  wire [22:0] prod_fraction__19;
  wire [7:0] incremented_sum__89;
  wire [27:0] wide_y__30;
  wire [7:0] x_bexpbs_difference__16;
  wire fraction_is_zero__31;
  wire [22:0] prod_fraction__92;
  wire [7:0] incremented_sum__107;
  wire [27:0] wide_y__63;
  wire [7:0] x_bexpbs_difference__31;
  wire fraction_is_zero__50;
  wire [22:0] prod_fraction__146;
  wire [7:0] incremented_sum__125;
  wire [27:0] wide_y__101;
  wire [7:0] x_bexpbs_difference__49;
  wire fraction_is_zero__69;
  wire [22:0] prod_fraction__200;
  wire [7:0] incremented_sum__143;
  wire [27:0] wide_y__139;
  wire [7:0] x_bexpbs_difference__67;
  wire [27:0] wide_y__13;
  wire [7:0] x_bexpbs_difference__7;
  wire [2:0] concat_167315;
  wire [7:0] x_bexp__126;
  wire [7:0] x_bexp__770;
  wire [27:0] wide_y__31;
  wire [7:0] sub_167321;
  wire [27:0] wide_y__64;
  wire [7:0] x_bexpbs_difference__32;
  wire [2:0] concat_167327;
  wire [7:0] x_bexp__251;
  wire [7:0] x_bexp__771;
  wire [27:0] wide_y__65;
  wire [7:0] sub_167333;
  wire [27:0] wide_y__102;
  wire [7:0] x_bexpbs_difference__50;
  wire [2:0] concat_167339;
  wire [7:0] x_bexp__395;
  wire [7:0] x_bexp__772;
  wire [27:0] wide_y__103;
  wire [7:0] sub_167345;
  wire [27:0] wide_y__140;
  wire [7:0] x_bexpbs_difference__68;
  wire [2:0] concat_167351;
  wire [7:0] x_bexp__539;
  wire [7:0] x_bexp__773;
  wire [27:0] wide_y__141;
  wire [7:0] sub_167357;
  wire [2:0] concat_167358;
  wire [7:0] x_bexp__54;
  wire [7:0] x_bexp__774;
  wire [27:0] wide_y__14;
  wire [7:0] sub_167364;
  wire result_sign__72;
  wire [22:0] x_fraction__126;
  wire [27:0] dropped__15;
  wire [2:0] concat_167372;
  wire [7:0] x_bexp__252;
  wire [7:0] x_bexp__775;
  wire [27:0] wide_y__66;
  wire [7:0] sub_167378;
  wire result_sign__152;
  wire [22:0] x_fraction__251;
  wire [27:0] dropped__32;
  wire [2:0] concat_167386;
  wire [7:0] x_bexp__396;
  wire [7:0] x_bexp__776;
  wire [27:0] wide_y__104;
  wire [7:0] sub_167392;
  wire result_sign__249;
  wire [22:0] x_fraction__395;
  wire [27:0] dropped__51;
  wire [2:0] concat_167400;
  wire [7:0] x_bexp__540;
  wire [7:0] x_bexp__777;
  wire [27:0] wide_y__142;
  wire [7:0] sub_167406;
  wire result_sign__346;
  wire [22:0] x_fraction__539;
  wire [27:0] dropped__70;
  wire result_sign__28;
  wire [22:0] x_fraction__54;
  wire [27:0] dropped__7;
  wire result_sign__73;
  wire [27:0] wide_x__30;
  wire result_sign__153;
  wire [22:0] x_fraction__252;
  wire [27:0] dropped__33;
  wire result_sign__154;
  wire [27:0] wide_x__63;
  wire x_sign__98;
  wire result_sign__250;
  wire [22:0] x_fraction__396;
  wire [27:0] dropped__52;
  wire nand_167448;
  wire result_sign__251;
  wire [27:0] wide_x__101;
  wire x_sign__134;
  wire result_sign__347;
  wire [22:0] x_fraction__540;
  wire [27:0] dropped__71;
  wire nand_167463;
  wire result_sign__348;
  wire [27:0] wide_x__139;
  wire result_sign__29;
  wire [27:0] wide_x__13;
  wire result_sign__76;
  wire result_sign__74;
  wire [27:0] wide_x__31;
  wire result_sign__155;
  wire [27:0] wide_x__64;
  wire result_sign__160;
  wire result_sign__156;
  wire [27:0] wide_x__65;
  wire result_sign__256;
  wire result_sign__252;
  wire [27:0] wide_x__102;
  wire result_sign__257;
  wire result_sign__253;
  wire [27:0] wide_x__103;
  wire result_sign__353;
  wire result_sign__349;
  wire [27:0] wide_x__140;
  wire result_sign__354;
  wire result_sign__350;
  wire [27:0] wide_x__141;
  wire result_sign__30;
  wire [27:0] wide_x__14;
  wire x_sign__32;
  wire prod_sign__15;
  wire [27:0] neg_167522;
  wire [27:0] sticky__47;
  wire result_sign__157;
  wire [27:0] wide_x__66;
  wire x_sign__63;
  wire prod_sign__31;
  wire [27:0] neg_167531;
  wire [27:0] sticky__100;
  wire result_sign__258;
  wire result_sign__254;
  wire [27:0] wide_x__104;
  wire x_sign__99;
  wire prod_sign__49;
  wire [27:0] neg_167541;
  wire [27:0] sticky__159;
  wire result_sign__355;
  wire result_sign__351;
  wire [27:0] wide_x__142;
  wire x_sign__135;
  wire prod_sign__67;
  wire [27:0] neg_167551;
  wire [27:0] sticky__218;
  wire x_sign__14;
  wire prod_sign__7;
  wire [27:0] neg_167556;
  wire [27:0] sticky__21;
  wire [27:0] xddend_y__15;
  wire x_sign__64;
  wire prod_sign__32;
  wire [27:0] neg_167565;
  wire [27:0] sticky__101;
  wire [27:0] xddend_y__31;
  wire x_sign__100;
  wire prod_sign__50;
  wire [27:0] neg_167574;
  wire [27:0] sticky__160;
  wire [27:0] xddend_y__49;
  wire x_sign__136;
  wire prod_sign__68;
  wire [27:0] neg_167583;
  wire [27:0] sticky__219;
  wire [27:0] xddend_y__67;
  wire [27:0] xddend_y__7;
  wire [24:0] sel_167594;
  wire result_sign__1050;
  wire [27:0] xddend_y__32;
  wire [24:0] sel_167601;
  wire result_sign__1051;
  wire [27:0] xddend_y__50;
  wire [24:0] sel_167608;
  wire result_sign__1052;
  wire [27:0] xddend_y__68;
  wire [24:0] sel_167615;
  wire result_sign__1053;
  wire [24:0] sel_167618;
  wire result_sign__1054;
  wire [24:0] sel_167623;
  wire result_sign__1055;
  wire [24:0] sel_167628;
  wire result_sign__1056;
  wire [24:0] sel_167633;
  wire result_sign__1057;
  wire [25:0] add_167640;
  wire [25:0] add_167643;
  wire [25:0] add_167646;
  wire [25:0] add_167649;
  wire [25:0] add_167650;
  wire [25:0] add_167653;
  wire [25:0] add_167656;
  wire [25:0] add_167659;
  wire [27:0] concat_167664;
  wire [27:0] concat_167667;
  wire [27:0] concat_167670;
  wire [27:0] concat_167673;
  wire [27:0] concat_167674;
  wire [27:0] concat_167677;
  wire [27:0] concat_167680;
  wire [27:0] concat_167683;
  wire [27:0] xbs_fraction__15;
  wire [27:0] xbs_fraction__31;
  wire [27:0] xbs_fraction__49;
  wire [27:0] xbs_fraction__67;
  wire [27:0] xbs_fraction__7;
  wire [27:0] reverse_167699;
  wire [27:0] xbs_fraction__32;
  wire [27:0] reverse_167701;
  wire [27:0] xbs_fraction__50;
  wire [27:0] reverse_167703;
  wire [27:0] xbs_fraction__68;
  wire [27:0] reverse_167705;
  wire [27:0] reverse_167706;
  wire [28:0] one_hot_167707;
  wire [27:0] reverse_167708;
  wire [28:0] one_hot_167709;
  wire [27:0] reverse_167710;
  wire [28:0] one_hot_167711;
  wire [27:0] reverse_167712;
  wire [28:0] one_hot_167713;
  wire [28:0] one_hot_167714;
  wire [4:0] encode_167715;
  wire [28:0] one_hot_167716;
  wire [4:0] encode_167717;
  wire [28:0] one_hot_167718;
  wire [4:0] encode_167719;
  wire [28:0] one_hot_167720;
  wire [4:0] encode_167721;
  wire [4:0] encode_167722;
  wire [4:0] encode_167724;
  wire [4:0] encode_167726;
  wire [4:0] encode_167728;
  wire cancel__16;
  wire carry_bit__15;
  wire [22:0] result_fraction__514;
  wire cancel__32;
  wire carry_bit__32;
  wire [22:0] result_fraction__581;
  wire cancel__51;
  wire carry_bit__51;
  wire [22:0] result_fraction__648;
  wire cancel__70;
  wire carry_bit__70;
  wire [22:0] result_fraction__723;
  wire cancel__7;
  wire carry_bit__7;
  wire [22:0] result_fraction__515;
  wire [27:0] leading_zeroes__15;
  wire cancel__33;
  wire carry_bit__33;
  wire [22:0] result_fraction__582;
  wire [27:0] leading_zeroes__32;
  wire cancel__52;
  wire carry_bit__52;
  wire [22:0] result_fraction__649;
  wire [27:0] leading_zeroes__51;
  wire cancel__71;
  wire carry_bit__71;
  wire [22:0] result_fraction__724;
  wire [27:0] leading_zeroes__70;
  wire [31:0] array_index_167783;
  wire [27:0] leading_zeroes__7;
  wire [26:0] carry_fraction__30;
  wire [27:0] add_167796;
  wire [27:0] leading_zeroes__33;
  wire [26:0] carry_fraction__63;
  wire [27:0] add_167809;
  wire [27:0] leading_zeroes__52;
  wire [26:0] carry_fraction__101;
  wire [27:0] add_167822;
  wire [27:0] leading_zeroes__71;
  wire [26:0] carry_fraction__139;
  wire [27:0] add_167835;
  wire [7:0] x_bexp__541;
  wire [26:0] carry_fraction__13;
  wire [27:0] add_167843;
  wire [2:0] concat_167844;
  wire [26:0] carry_fraction__31;
  wire [26:0] cancel_fraction__15;
  wire [26:0] carry_fraction__64;
  wire [27:0] add_167853;
  wire [2:0] concat_167854;
  wire [26:0] carry_fraction__65;
  wire [26:0] cancel_fraction__32;
  wire [26:0] carry_fraction__102;
  wire [27:0] add_167863;
  wire [2:0] concat_167864;
  wire [26:0] carry_fraction__103;
  wire [26:0] cancel_fraction__51;
  wire result_sign__1058;
  wire [26:0] carry_fraction__140;
  wire [27:0] add_167875;
  wire [2:0] concat_167876;
  wire [26:0] carry_fraction__141;
  wire [26:0] cancel_fraction__70;
  wire result_sign__1059;
  wire [2:0] concat_167881;
  wire [26:0] carry_fraction__14;
  wire [26:0] cancel_fraction__7;
  wire [26:0] shifted_fraction__15;
  wire [2:0] concat_167885;
  wire [26:0] carry_fraction__66;
  wire [26:0] cancel_fraction__33;
  wire [26:0] shifted_fraction__32;
  wire [2:0] concat_167889;
  wire [26:0] carry_fraction__104;
  wire [26:0] cancel_fraction__52;
  wire [26:0] shifted_fraction__51;
  wire [2:0] concat_167895;
  wire [26:0] carry_fraction__142;
  wire [26:0] cancel_fraction__71;
  wire [26:0] shifted_fraction__70;
  wire [26:0] shifted_fraction__7;
  wire result_sign__1060;
  wire [26:0] shifted_fraction__33;
  wire result_sign__1061;
  wire [26:0] shifted_fraction__52;
  wire result_sign__1062;
  wire result_sign__1111;
  wire [1:0] add_167911;
  wire [26:0] shifted_fraction__71;
  wire result_sign__1063;
  wire result_sign__1115;
  wire [1:0] add_167917;
  wire [7:0] x_bexp__778;
  wire result_sign__747;
  wire [22:0] x_fraction__541;
  wire result_sign__1064;
  wire [2:0] normal_chunk__15;
  wire [2:0] fraction_shift__249;
  wire [1:0] half_way_chunk__15;
  wire result_sign__1065;
  wire [2:0] normal_chunk__32;
  wire [2:0] fraction_shift__284;
  wire [1:0] half_way_chunk__32;
  wire result_sign__1066;
  wire [2:0] normal_chunk__51;
  wire [2:0] fraction_shift__319;
  wire [1:0] half_way_chunk__51;
  wire result_sign__1067;
  wire [2:0] normal_chunk__70;
  wire [2:0] fraction_shift__354;
  wire [1:0] half_way_chunk__70;
  wire ne_167958;
  wire [2:0] normal_chunk__7;
  wire [2:0] fraction_shift__250;
  wire [1:0] half_way_chunk__7;
  wire result_sign__442;
  wire [24:0] add_167970;
  wire [2:0] normal_chunk__33;
  wire [2:0] fraction_shift__285;
  wire [1:0] half_way_chunk__33;
  wire result_sign__539;
  wire [24:0] add_167980;
  wire [2:0] normal_chunk__52;
  wire [2:0] fraction_shift__320;
  wire [1:0] half_way_chunk__52;
  wire result_sign__639;
  wire [24:0] add_167990;
  wire [9:0] exp__221;
  wire [2:0] normal_chunk__71;
  wire [2:0] fraction_shift__355;
  wire [1:0] half_way_chunk__71;
  wire result_sign__749;
  wire [24:0] add_168001;
  wire [9:0] exp__303;
  wire [9:0] sign_ext_168003;
  wire [23:0] x_fraction__543;
  wire result_sign__443;
  wire [24:0] add_168009;
  wire do_round_up__31;
  wire result_sign__540;
  wire [24:0] add_168016;
  wire do_round_up__66;
  wire result_sign__640;
  wire [24:0] add_168023;
  wire do_round_up__105;
  wire [9:0] exp__223;
  wire result_sign__750;
  wire [24:0] add_168032;
  wire do_round_up__144;
  wire [9:0] exp__305;
  wire [23:0] x_fraction__545;
  wire result_sign__824;
  wire result_sign__825;
  wire do_round_up__14;
  wire [27:0] rounded_fraction__15;
  wire do_round_up__67;
  wire [27:0] rounded_fraction__32;
  wire do_round_up__106;
  wire [27:0] rounded_fraction__51;
  wire do_round_up__145;
  wire [27:0] rounded_fraction__70;
  wire [24:0] concat_168059;
  wire [24:0] concat_168060;
  wire [27:0] rounded_fraction__7;
  wire result_sign__444;
  wire [7:0] x_bexp__586;
  wire rounding_carry__15;
  wire [27:0] rounded_fraction__33;
  wire result_sign__541;
  wire [7:0] x_bexp__604;
  wire rounding_carry__32;
  wire [27:0] rounded_fraction__52;
  wire result_sign__641;
  wire [7:0] x_bexp__622;
  wire rounding_carry__51;
  wire [24:0] sel_168073;
  wire [27:0] rounded_fraction__71;
  wire result_sign__751;
  wire [7:0] x_bexp__640;
  wire rounding_carry__70;
  wire [24:0] sel_168078;
  wire result_sign__445;
  wire [7:0] x_bexp__587;
  wire rounding_carry__7;
  wire result_sign__542;
  wire [7:0] x_bexp__605;
  wire rounding_carry__33;
  wire result_sign__642;
  wire [7:0] x_bexp__623;
  wire rounding_carry__52;
  wire result_sign__946;
  wire [22:0] fraction__495;
  wire result_sign__752;
  wire [7:0] x_bexp__641;
  wire rounding_carry__71;
  wire result_sign__954;
  wire [22:0] fraction__674;
  wire result_sign__446;
  wire [8:0] add_168106;
  wire result_sign__543;
  wire [8:0] add_168112;
  wire result_sign__643;
  wire [8:0] add_168118;
  wire [23:0] fraction__497;
  wire result_sign__753;
  wire [8:0] add_168128;
  wire [23:0] fraction__676;
  wire result_sign__447;
  wire [8:0] add_168136;
  wire result_sign__544;
  wire [8:0] add_168145;
  wire result_sign__644;
  wire [8:0] add_168154;
  wire do_round_up__107;
  wire [23:0] add_168163;
  wire result_sign__754;
  wire [8:0] add_168165;
  wire do_round_up__146;
  wire [23:0] add_168174;
  wire [9:0] add_168180;
  wire [9:0] add_168188;
  wire [9:0] add_168196;
  wire [23:0] fraction__499;
  wire [9:0] add_168206;
  wire [23:0] fraction__678;
  wire [9:0] add_168211;
  wire [9:0] wide_exponent__45;
  wire [9:0] add_168216;
  wire [9:0] wide_exponent__94;
  wire [9:0] add_168221;
  wire [9:0] wide_exponent__151;
  wire [9:0] add_168227;
  wire [9:0] add_168228;
  wire [9:0] wide_exponent__208;
  wire [9:0] add_168234;
  wire [9:0] wide_exponent__19;
  wire [9:0] wide_exponent__46;
  wire [9:0] wide_exponent__95;
  wire [9:0] wide_exponent__96;
  wire [9:0] wide_exponent__152;
  wire [9:0] wide_exponent__153;
  wire [9:0] exp__227;
  wire [9:0] wide_exponent__209;
  wire [9:0] wide_exponent__210;
  wire [9:0] exp__309;
  wire [9:0] wide_exponent__20;
  wire [7:0] high_exp__375;
  wire [22:0] result_fraction__781;
  wire [7:0] high_exp__376;
  wire [22:0] result_fraction__782;
  wire [7:0] high_exp__117;
  wire [22:0] result_fraction__516;
  wire [7:0] high_exp__118;
  wire [22:0] result_fraction__517;
  wire [9:0] wide_exponent__97;
  wire [7:0] high_exp__407;
  wire [22:0] result_fraction__814;
  wire [7:0] high_exp__408;
  wire [22:0] result_fraction__815;
  wire [7:0] high_exp__182;
  wire [22:0] result_fraction__583;
  wire [7:0] high_exp__183;
  wire [22:0] result_fraction__584;
  wire [9:0] wide_exponent__154;
  wire [7:0] high_exp__439;
  wire [22:0] result_fraction__847;
  wire [7:0] high_exp__440;
  wire [22:0] result_fraction__848;
  wire [7:0] high_exp__249;
  wire [22:0] result_fraction__650;
  wire [7:0] high_exp__250;
  wire [22:0] result_fraction__651;
  wire [9:0] wide_exponent__211;
  wire [7:0] high_exp__471;
  wire [22:0] result_fraction__880;
  wire [7:0] high_exp__472;
  wire [22:0] result_fraction__881;
  wire [7:0] high_exp__321;
  wire [22:0] result_fraction__725;
  wire [7:0] high_exp__322;
  wire [22:0] result_fraction__726;
  wire [7:0] high_exp__361;
  wire [22:0] result_fraction__766;
  wire [7:0] high_exp__362;
  wire [22:0] result_fraction__767;
  wire [7:0] high_exp__119;
  wire [22:0] result_fraction__518;
  wire [7:0] high_exp__120;
  wire [22:0] result_fraction__519;
  wire ne_168304;
  wire ne_168306;
  wire eq_168307;
  wire eq_168308;
  wire eq_168309;
  wire eq_168310;
  wire [7:0] high_exp__393;
  wire [22:0] result_fraction__799;
  wire [7:0] high_exp__394;
  wire [22:0] result_fraction__800;
  wire [7:0] high_exp__184;
  wire [22:0] result_fraction__585;
  wire [7:0] high_exp__185;
  wire [22:0] result_fraction__586;
  wire ne_168322;
  wire ne_168324;
  wire eq_168325;
  wire eq_168326;
  wire eq_168327;
  wire eq_168328;
  wire [7:0] high_exp__425;
  wire [22:0] result_fraction__832;
  wire [7:0] high_exp__426;
  wire [22:0] result_fraction__833;
  wire [7:0] high_exp__251;
  wire [22:0] result_fraction__652;
  wire [7:0] high_exp__252;
  wire [22:0] result_fraction__653;
  wire ne_168340;
  wire ne_168342;
  wire eq_168343;
  wire eq_168344;
  wire eq_168345;
  wire eq_168346;
  wire [8:0] result_exp__163;
  wire [7:0] high_exp__457;
  wire [22:0] result_fraction__865;
  wire [7:0] high_exp__458;
  wire [22:0] result_fraction__866;
  wire [7:0] high_exp__323;
  wire [22:0] result_fraction__727;
  wire [7:0] high_exp__324;
  wire [22:0] result_fraction__728;
  wire ne_168360;
  wire ne_168362;
  wire eq_168363;
  wire eq_168364;
  wire eq_168365;
  wire eq_168366;
  wire [8:0] result_exp__223;
  wire ne_168371;
  wire ne_168373;
  wire eq_168374;
  wire eq_168375;
  wire eq_168376;
  wire eq_168377;
  wire ne_168386;
  wire ne_168388;
  wire eq_168389;
  wire eq_168390;
  wire eq_168391;
  wire eq_168392;
  wire ne_168401;
  wire ne_168403;
  wire eq_168404;
  wire eq_168405;
  wire eq_168406;
  wire eq_168407;
  wire [8:0] result_exp__165;
  wire ne_168417;
  wire ne_168419;
  wire eq_168420;
  wire eq_168421;
  wire eq_168422;
  wire eq_168423;
  wire [7:0] high_exp__326;
  wire [22:0] result_fraction__730;
  wire [22:0] result_fraction__729;
  wire [8:0] result_exp__225;
  wire [8:0] wide_exponent__47;
  wire has_pos_inf__15;
  wire has_neg_inf__15;
  wire [8:0] wide_exponent__98;
  wire has_pos_inf__32;
  wire has_neg_inf__32;
  wire [8:0] wide_exponent__155;
  wire has_pos_inf__51;
  wire has_neg_inf__51;
  wire [8:0] wide_exponent__212;
  wire has_pos_inf__70;
  wire has_neg_inf__70;
  wire is_result_nan__147;
  wire ne_168472;
  wire [8:0] wide_exponent__21;
  wire has_pos_inf__7;
  wire has_neg_inf__7;
  wire [8:0] wide_exponent__99;
  wire has_pos_inf__33;
  wire has_neg_inf__33;
  wire [8:0] wide_exponent__156;
  wire has_pos_inf__52;
  wire has_neg_inf__52;
  wire and_reduce_168506;
  wire [8:0] wide_exponent__213;
  wire has_pos_inf__71;
  wire has_neg_inf__71;
  wire is_result_nan__146;
  wire has_inf_arg__76;
  wire and_reduce_168520;
  wire is_result_nan__31;
  wire is_operand_inf__15;
  wire and_reduce_168533;
  wire is_result_nan__66;
  wire is_operand_inf__32;
  wire and_reduce_168546;
  wire is_result_nan__105;
  wire is_operand_inf__51;
  wire and_reduce_168560;
  wire [7:0] high_exp__255;
  wire is_result_nan__144;
  wire is_operand_inf__70;
  wire and_reduce_168576;
  wire [7:0] high_exp__328;
  wire is_result_nan__14;
  wire is_operand_inf__7;
  wire and_reduce_168584;
  wire [2:0] fraction_shift__378;
  wire [2:0] fraction_shift__251;
  wire [7:0] high_exp__121;
  wire is_result_nan__67;
  wire is_operand_inf__33;
  wire and_reduce_168595;
  wire [2:0] fraction_shift__396;
  wire [2:0] fraction_shift__286;
  wire [7:0] high_exp__186;
  wire is_result_nan__106;
  wire is_operand_inf__52;
  wire and_reduce_168606;
  wire [2:0] fraction_shift__414;
  wire [2:0] fraction_shift__321;
  wire is_subnormal__55;
  wire [7:0] high_exp__253;
  wire [7:0] result_exp__167;
  wire is_result_nan__145;
  wire is_operand_inf__71;
  wire and_reduce_168619;
  wire [2:0] fraction_shift__432;
  wire [2:0] fraction_shift__356;
  wire is_subnormal__75;
  wire [7:0] high_exp__325;
  wire [7:0] result_exp__227;
  wire [2:0] fraction_shift__379;
  wire [2:0] fraction_shift__252;
  wire [7:0] high_exp__122;
  wire [2:0] fraction_shift__48;
  wire result_sign__448;
  wire [7:0] result_exponent__16;
  wire [2:0] fraction_shift__397;
  wire [2:0] fraction_shift__287;
  wire [7:0] high_exp__187;
  wire [2:0] fraction_shift__98;
  wire result_sign__545;
  wire [7:0] result_exponent__32;
  wire [2:0] fraction_shift__415;
  wire [2:0] fraction_shift__322;
  wire [7:0] high_exp__254;
  wire [7:0] result_exp__168;
  wire [2:0] fraction_shift__155;
  wire result_sign__645;
  wire [7:0] result_exponent__51;
  wire result_sign__646;
  wire [2:0] fraction_shift__433;
  wire [2:0] fraction_shift__357;
  wire [7:0] high_exp__327;
  wire [7:0] result_exp__228;
  wire [2:0] fraction_shift__212;
  wire result_sign__755;
  wire [7:0] result_exponent__70;
  wire result_sign__756;
  wire [2:0] fraction_shift__21;
  wire result_sign__449;
  wire [7:0] result_exponent__7;
  wire [27:0] shrl_168675;
  wire [2:0] fraction_shift__99;
  wire result_sign__546;
  wire [7:0] result_exponent__33;
  wire [27:0] shrl_168682;
  wire [2:0] fraction_shift__156;
  wire result_sign__647;
  wire [7:0] result_exponent__52;
  wire result_sign__648;
  wire [27:0] shrl_168691;
  wire [2:0] fraction_shift__213;
  wire result_sign__757;
  wire [7:0] result_exponent__71;
  wire result_sign__758;
  wire [27:0] shrl_168702;
  wire [27:0] shrl_168707;
  wire [22:0] result_fraction__93;
  wire [8:0] sum__16;
  wire [27:0] shrl_168713;
  wire [22:0] result_fraction__196;
  wire [8:0] sum__34;
  wire [27:0] shrl_168719;
  wire [22:0] result_fraction__313;
  wire [22:0] result_fraction__319;
  wire [8:0] sum__53;
  wire [27:0] shrl_168728;
  wire [22:0] result_fraction__430;
  wire [22:0] result_fraction__436;
  wire [8:0] sum__72;
  wire [22:0] result_fraction__40;
  wire [8:0] sum__8;
  wire [22:0] result_fraction__94;
  wire [22:0] nan_fraction__96;
  wire [22:0] result_fraction__197;
  wire [8:0] sum__35;
  wire [22:0] result_fraction__198;
  wire [22:0] nan_fraction__123;
  wire [22:0] result_fraction__314;
  wire [8:0] sum__54;
  wire [22:0] result_fraction__315;
  wire [22:0] nan_fraction__151;
  wire [22:0] result_fraction__321;
  wire [22:0] nan_fraction__153;
  wire [22:0] result_fraction__431;
  wire [8:0] sum__73;
  wire [22:0] result_fraction__432;
  wire [22:0] nan_fraction__180;
  wire [22:0] result_fraction__438;
  wire [22:0] nan_fraction__182;
  wire [22:0] result_fraction__41;
  wire [22:0] nan_fraction__97;
  wire [22:0] result_fraction__95;
  wire [7:0] prod_bexp__66;
  wire [7:0] x_bexp__779;
  wire [22:0] result_fraction__199;
  wire [22:0] nan_fraction__124;
  wire [22:0] result_fraction__200;
  wire [7:0] prod_bexp__131;
  wire [7:0] x_bexp__780;
  wire [22:0] result_fraction__316;
  wire [22:0] nan_fraction__152;
  wire [22:0] result_fraction__317;
  wire [22:0] result_fraction__323;
  wire [7:0] prod_bexp__203;
  wire [7:0] x_bexp__781;
  wire [22:0] result_fraction__433;
  wire [22:0] nan_fraction__181;
  wire [22:0] result_fraction__434;
  wire [22:0] result_fraction__440;
  wire [7:0] prod_bexp__275;
  wire [7:0] x_bexp__782;
  wire [22:0] result_fraction__42;
  wire [7:0] prod_bexp__30;
  wire [7:0] x_bexp__783;
  wire fraction_is_zero__15;
  wire [22:0] prod_fraction__48;
  wire [7:0] incremented_sum__90;
  wire [22:0] result_fraction__201;
  wire [7:0] prod_bexp__132;
  wire [7:0] x_bexp__784;
  wire fraction_is_zero__32;
  wire [22:0] prod_fraction__97;
  wire [7:0] incremented_sum__108;
  wire [22:0] result_fraction__318;
  wire [22:0] result_fraction__479;
  wire [7:0] prod_bexp__204;
  wire [7:0] x_bexp__785;
  wire fraction_is_zero__51;
  wire [22:0] prod_fraction__151;
  wire [7:0] incremented_sum__126;
  wire [22:0] result_fraction__435;
  wire [22:0] result_fraction__480;
  wire [7:0] prod_bexp__276;
  wire [7:0] x_bexp__786;
  wire fraction_is_zero__70;
  wire [22:0] prod_fraction__205;
  wire [7:0] incremented_sum__144;
  wire fraction_is_zero__7;
  wire [22:0] prod_fraction__22;
  wire [7:0] incremented_sum__91;
  wire [27:0] wide_y__32;
  wire [7:0] x_bexpbs_difference__17;
  wire fraction_is_zero__33;
  wire [22:0] prod_fraction__98;
  wire [7:0] incremented_sum__109;
  wire [27:0] wide_y__67;
  wire [7:0] x_bexpbs_difference__33;
  wire fraction_is_zero__52;
  wire [22:0] prod_fraction__152;
  wire [7:0] incremented_sum__127;
  wire [27:0] wide_y__105;
  wire [7:0] x_bexpbs_difference__51;
  wire fraction_is_zero__71;
  wire [22:0] prod_fraction__206;
  wire [7:0] incremented_sum__145;
  wire [27:0] wide_y__143;
  wire [7:0] x_bexpbs_difference__69;
  wire [27:0] wide_y__15;
  wire [7:0] x_bexpbs_difference__8;
  wire [2:0] concat_168936;
  wire [7:0] x_bexp__134;
  wire [7:0] x_bexp__787;
  wire [27:0] wide_y__33;
  wire [7:0] sub_168942;
  wire [27:0] wide_y__68;
  wire [7:0] x_bexpbs_difference__34;
  wire [2:0] concat_168948;
  wire [7:0] x_bexp__267;
  wire [7:0] x_bexp__788;
  wire [27:0] wide_y__69;
  wire [7:0] sub_168954;
  wire [27:0] wide_y__106;
  wire [7:0] x_bexpbs_difference__52;
  wire [2:0] concat_168960;
  wire [7:0] x_bexp__411;
  wire [7:0] x_bexp__789;
  wire [27:0] wide_y__107;
  wire [7:0] sub_168966;
  wire [27:0] wide_y__144;
  wire [7:0] x_bexpbs_difference__70;
  wire [2:0] concat_168972;
  wire [7:0] x_bexp__555;
  wire [7:0] x_bexp__790;
  wire [27:0] wide_y__145;
  wire [7:0] sub_168978;
  wire [2:0] concat_168979;
  wire [7:0] x_bexp__62;
  wire [7:0] x_bexp__791;
  wire [27:0] wide_y__16;
  wire [7:0] sub_168985;
  wire result_sign__77;
  wire [22:0] x_fraction__134;
  wire [27:0] dropped__16;
  wire [2:0] concat_168993;
  wire [7:0] x_bexp__268;
  wire [7:0] x_bexp__792;
  wire [27:0] wide_y__70;
  wire [7:0] sub_168999;
  wire result_sign__162;
  wire [22:0] x_fraction__267;
  wire [27:0] dropped__34;
  wire [2:0] concat_169007;
  wire [7:0] x_bexp__412;
  wire [7:0] x_bexp__793;
  wire [27:0] wide_y__108;
  wire [7:0] sub_169013;
  wire result_sign__259;
  wire [22:0] x_fraction__411;
  wire [27:0] dropped__53;
  wire [2:0] concat_169021;
  wire [7:0] x_bexp__556;
  wire [7:0] x_bexp__794;
  wire [27:0] wide_y__146;
  wire [7:0] sub_169027;
  wire result_sign__356;
  wire [22:0] x_fraction__555;
  wire [27:0] dropped__72;
  wire result_sign__33;
  wire [22:0] x_fraction__62;
  wire [27:0] dropped__8;
  wire result_sign__78;
  wire [27:0] wide_x__32;
  wire result_sign__163;
  wire [22:0] x_fraction__268;
  wire [27:0] dropped__35;
  wire result_sign__164;
  wire [27:0] wide_x__67;
  wire [7:0] high_exp__485;
  wire result_sign__260;
  wire [22:0] x_fraction__412;
  wire [27:0] dropped__54;
  wire result_sign__261;
  wire [27:0] wide_x__105;
  wire [7:0] high_exp__490;
  wire result_sign__357;
  wire [22:0] x_fraction__556;
  wire [27:0] dropped__73;
  wire x_sign__137;
  wire result_sign__358;
  wire [27:0] wide_x__143;
  wire result_sign__34;
  wire [27:0] wide_x__15;
  wire result_sign__79;
  wire [27:0] wide_x__33;
  wire result_sign__165;
  wire [27:0] wide_x__68;
  wire result_sign__166;
  wire [27:0] wide_x__69;
  wire result_sign__262;
  wire [27:0] wide_x__106;
  wire result_sign__263;
  wire [27:0] wide_x__107;
  wire result_sign__359;
  wire [27:0] wide_x__144;
  wire result_sign__364;
  wire result_sign__360;
  wire [27:0] wide_x__145;
  wire result_sign__35;
  wire [27:0] wide_x__16;
  wire x_sign__34;
  wire prod_sign__16;
  wire [27:0] neg_169140;
  wire [27:0] sticky__50;
  wire result_sign__167;
  wire [27:0] wide_x__70;
  wire x_sign__67;
  wire prod_sign__33;
  wire [27:0] neg_169149;
  wire [27:0] sticky__106;
  wire result_sign__268;
  wire result_sign__264;
  wire [27:0] wide_x__108;
  wire x_sign__103;
  wire prod_sign__51;
  wire [27:0] neg_169159;
  wire [27:0] sticky__165;
  wire result_sign__365;
  wire result_sign__361;
  wire [27:0] wide_x__146;
  wire x_sign__139;
  wire prod_sign__69;
  wire [27:0] neg_169169;
  wire [27:0] sticky__224;
  wire x_sign__16;
  wire prod_sign__8;
  wire [27:0] neg_169174;
  wire [27:0] sticky__24;
  wire [27:0] xddend_y__16;
  wire x_sign__68;
  wire prod_sign__34;
  wire [27:0] neg_169183;
  wire [27:0] sticky__107;
  wire [27:0] xddend_y__33;
  wire x_sign__104;
  wire prod_sign__52;
  wire [27:0] neg_169192;
  wire [27:0] sticky__166;
  wire [27:0] xddend_y__51;
  wire x_sign__140;
  wire prod_sign__70;
  wire [27:0] neg_169201;
  wire [27:0] sticky__225;
  wire [27:0] xddend_y__69;
  wire [27:0] xddend_y__8;
  wire [24:0] sel_169212;
  wire result_sign__1068;
  wire [27:0] xddend_y__34;
  wire [24:0] sel_169219;
  wire result_sign__1069;
  wire [27:0] xddend_y__52;
  wire [24:0] sel_169226;
  wire result_sign__1070;
  wire [27:0] xddend_y__70;
  wire [24:0] sel_169233;
  wire result_sign__1071;
  wire [24:0] sel_169236;
  wire result_sign__1072;
  wire [24:0] sel_169241;
  wire result_sign__1073;
  wire [24:0] sel_169246;
  wire result_sign__1074;
  wire [24:0] sel_169251;
  wire result_sign__1075;
  wire [25:0] add_169258;
  wire [25:0] add_169261;
  wire [25:0] add_169264;
  wire [25:0] add_169267;
  wire [25:0] add_169268;
  wire [25:0] add_169271;
  wire [25:0] add_169274;
  wire [25:0] add_169277;
  wire [27:0] concat_169282;
  wire [27:0] concat_169285;
  wire [27:0] concat_169288;
  wire [27:0] concat_169291;
  wire [27:0] concat_169292;
  wire [27:0] concat_169295;
  wire [27:0] concat_169298;
  wire [27:0] concat_169301;
  wire [27:0] xbs_fraction__16;
  wire [27:0] xbs_fraction__33;
  wire [27:0] xbs_fraction__51;
  wire [27:0] xbs_fraction__69;
  wire [27:0] xbs_fraction__8;
  wire [27:0] reverse_169317;
  wire [27:0] xbs_fraction__34;
  wire [27:0] reverse_169319;
  wire [27:0] xbs_fraction__52;
  wire [27:0] reverse_169321;
  wire [27:0] xbs_fraction__70;
  wire [27:0] reverse_169323;
  wire [27:0] reverse_169324;
  wire [28:0] one_hot_169325;
  wire [27:0] reverse_169326;
  wire [28:0] one_hot_169327;
  wire [27:0] reverse_169328;
  wire [28:0] one_hot_169329;
  wire [27:0] reverse_169330;
  wire [28:0] one_hot_169331;
  wire [28:0] one_hot_169332;
  wire [4:0] encode_169333;
  wire [28:0] one_hot_169334;
  wire [4:0] encode_169335;
  wire [28:0] one_hot_169336;
  wire [4:0] encode_169337;
  wire [28:0] one_hot_169338;
  wire [4:0] encode_169339;
  wire [4:0] encode_169340;
  wire [4:0] encode_169342;
  wire [4:0] encode_169344;
  wire [4:0] encode_169346;
  wire cancel__17;
  wire carry_bit__16;
  wire [22:0] result_fraction__520;
  wire cancel__34;
  wire carry_bit__34;
  wire [22:0] result_fraction__587;
  wire cancel__53;
  wire carry_bit__53;
  wire [22:0] result_fraction__654;
  wire cancel__72;
  wire carry_bit__72;
  wire [22:0] result_fraction__731;
  wire cancel__8;
  wire carry_bit__8;
  wire [22:0] result_fraction__521;
  wire [27:0] leading_zeroes__16;
  wire cancel__35;
  wire carry_bit__35;
  wire [22:0] result_fraction__588;
  wire [27:0] leading_zeroes__34;
  wire cancel__54;
  wire carry_bit__54;
  wire [22:0] result_fraction__655;
  wire [27:0] leading_zeroes__53;
  wire cancel__73;
  wire carry_bit__73;
  wire [22:0] result_fraction__732;
  wire [27:0] leading_zeroes__72;
  wire [27:0] leading_zeroes__8;
  wire [26:0] carry_fraction__32;
  wire [27:0] add_169413;
  wire [27:0] leading_zeroes__35;
  wire [26:0] carry_fraction__67;
  wire [27:0] add_169426;
  wire [27:0] leading_zeroes__54;
  wire [26:0] carry_fraction__105;
  wire [27:0] add_169439;
  wire [27:0] leading_zeroes__73;
  wire [26:0] carry_fraction__143;
  wire [27:0] add_169452;
  wire [31:0] array_index_169453;
  wire [26:0] carry_fraction__15;
  wire [27:0] add_169460;
  wire [2:0] concat_169461;
  wire [26:0] carry_fraction__33;
  wire [26:0] cancel_fraction__16;
  wire result_sign__617;
  wire [26:0] carry_fraction__68;
  wire [27:0] add_169471;
  wire [2:0] concat_169472;
  wire [26:0] carry_fraction__69;
  wire [26:0] cancel_fraction__34;
  wire result_sign__724;
  wire [26:0] carry_fraction__106;
  wire [27:0] add_169482;
  wire [2:0] concat_169483;
  wire [26:0] carry_fraction__107;
  wire [26:0] cancel_fraction__53;
  wire result_sign__748;
  wire [26:0] carry_fraction__144;
  wire [27:0] add_169493;
  wire [2:0] concat_169494;
  wire [26:0] carry_fraction__145;
  wire [26:0] cancel_fraction__72;
  wire result_sign__760;
  wire [7:0] x_bexp__557;
  wire [2:0] concat_169499;
  wire [26:0] carry_fraction__16;
  wire [26:0] cancel_fraction__8;
  wire [26:0] shifted_fraction__16;
  wire [2:0] concat_169505;
  wire [26:0] carry_fraction__70;
  wire [26:0] cancel_fraction__35;
  wire [26:0] shifted_fraction__34;
  wire [2:0] concat_169511;
  wire [26:0] carry_fraction__108;
  wire [26:0] cancel_fraction__54;
  wire [26:0] shifted_fraction__53;
  wire [2:0] concat_169517;
  wire [26:0] carry_fraction__146;
  wire [26:0] cancel_fraction__73;
  wire [26:0] shifted_fraction__72;
  wire [26:0] shifted_fraction__8;
  wire result_sign__1076;
  wire result_sign__452;
  wire [8:0] add_169527;
  wire [26:0] shifted_fraction__35;
  wire result_sign__1077;
  wire result_sign__549;
  wire [8:0] add_169532;
  wire [26:0] shifted_fraction__54;
  wire result_sign__1078;
  wire result_sign__651;
  wire [8:0] add_169537;
  wire [26:0] shifted_fraction__73;
  wire result_sign__1079;
  wire result_sign__763;
  wire [8:0] add_169542;
  wire [7:0] x_bexp__795;
  wire result_sign__759;
  wire [22:0] x_fraction__557;
  wire result_sign__1080;
  wire [2:0] normal_chunk__16;
  wire [2:0] fraction_shift__253;
  wire [1:0] half_way_chunk__16;
  wire result_sign__1081;
  wire [2:0] normal_chunk__34;
  wire [2:0] fraction_shift__288;
  wire [1:0] half_way_chunk__34;
  wire result_sign__1082;
  wire [2:0] normal_chunk__53;
  wire [2:0] fraction_shift__323;
  wire [1:0] half_way_chunk__53;
  wire result_sign__1083;
  wire [2:0] normal_chunk__72;
  wire [2:0] fraction_shift__358;
  wire [1:0] half_way_chunk__72;
  wire ne_169586;
  wire [2:0] normal_chunk__8;
  wire [2:0] fraction_shift__254;
  wire [1:0] half_way_chunk__8;
  wire result_sign__450;
  wire [24:0] add_169598;
  wire [9:0] exp__68;
  wire [2:0] normal_chunk__35;
  wire [2:0] fraction_shift__289;
  wire [1:0] half_way_chunk__35;
  wire result_sign__547;
  wire [24:0] add_169609;
  wire [9:0] exp__147;
  wire [2:0] normal_chunk__54;
  wire [2:0] fraction_shift__324;
  wire [1:0] half_way_chunk__54;
  wire result_sign__649;
  wire [24:0] add_169620;
  wire [9:0] exp__229;
  wire [2:0] normal_chunk__73;
  wire [2:0] fraction_shift__359;
  wire [1:0] half_way_chunk__73;
  wire result_sign__761;
  wire [24:0] add_169631;
  wire [9:0] exp__311;
  wire [23:0] x_fraction__559;
  wire result_sign__451;
  wire [24:0] add_169639;
  wire do_round_up__33;
  wire [9:0] exp__69;
  wire result_sign__548;
  wire [24:0] add_169648;
  wire do_round_up__70;
  wire [9:0] exp__149;
  wire result_sign__650;
  wire [24:0] add_169657;
  wire do_round_up__109;
  wire [9:0] exp__231;
  wire result_sign__762;
  wire [24:0] add_169666;
  wire do_round_up__148;
  wire [9:0] exp__313;
  wire [23:0] x_fraction__561;
  wire result_sign__826;
  wire result_sign__827;
  wire do_round_up__16;
  wire [27:0] rounded_fraction__16;
  wire do_round_up__71;
  wire [27:0] rounded_fraction__34;
  wire do_round_up__110;
  wire [27:0] rounded_fraction__53;
  wire do_round_up__149;
  wire [27:0] rounded_fraction__72;
  wire [27:0] rounded_fraction__8;
  wire result_sign__453;
  wire [7:0] x_bexp__588;
  wire rounding_carry__16;
  wire [24:0] sel_169701;
  wire [27:0] rounded_fraction__35;
  wire result_sign__550;
  wire [7:0] x_bexp__606;
  wire rounding_carry__34;
  wire [24:0] sel_169706;
  wire [27:0] rounded_fraction__54;
  wire result_sign__652;
  wire [7:0] x_bexp__624;
  wire rounding_carry__53;
  wire [24:0] sel_169711;
  wire [27:0] rounded_fraction__73;
  wire result_sign__764;
  wire [7:0] x_bexp__642;
  wire rounding_carry__72;
  wire [24:0] sel_169716;
  wire result_sign__454;
  wire [7:0] x_bexp__589;
  wire rounding_carry__8;
  wire result_sign__933;
  wire [22:0] fraction__158;
  wire result_sign__551;
  wire [7:0] x_bexp__607;
  wire rounding_carry__35;
  wire result_sign__939;
  wire [22:0] fraction__334;
  wire result_sign__653;
  wire [7:0] x_bexp__625;
  wire rounding_carry__54;
  wire result_sign__947;
  wire [22:0] fraction__513;
  wire result_sign__765;
  wire [7:0] x_bexp__643;
  wire rounding_carry__73;
  wire result_sign__955;
  wire [22:0] fraction__692;
  wire result_sign__455;
  wire [8:0] add_169748;
  wire [23:0] fraction__159;
  wire result_sign__552;
  wire [8:0] add_169758;
  wire [23:0] fraction__336;
  wire result_sign__654;
  wire [8:0] add_169768;
  wire [23:0] fraction__515;
  wire result_sign__766;
  wire [8:0] add_169778;
  wire [23:0] fraction__694;
  wire result_sign__456;
  wire [8:0] add_169786;
  wire do_round_up__34;
  wire [23:0] add_169795;
  wire result_sign__553;
  wire [8:0] add_169797;
  wire do_round_up__72;
  wire [23:0] add_169806;
  wire result_sign__655;
  wire [8:0] add_169808;
  wire do_round_up__111;
  wire [23:0] add_169817;
  wire result_sign__767;
  wire [8:0] add_169819;
  wire do_round_up__150;
  wire [23:0] add_169828;
  wire [9:0] add_169834;
  wire [23:0] fraction__160;
  wire [9:0] add_169844;
  wire [23:0] fraction__338;
  wire [9:0] add_169854;
  wire [23:0] fraction__517;
  wire [9:0] add_169864;
  wire [23:0] fraction__696;
  wire [9:0] add_169869;
  wire [9:0] wide_exponent__48;
  wire [9:0] add_169875;
  wire [9:0] add_169876;
  wire [9:0] wide_exponent__100;
  wire [9:0] add_169882;
  wire [9:0] add_169883;
  wire [9:0] wide_exponent__157;
  wire [9:0] add_169889;
  wire [9:0] add_169890;
  wire [9:0] wide_exponent__214;
  wire [9:0] add_169896;
  wire [9:0] wide_exponent__22;
  wire [9:0] wide_exponent__49;
  wire [9:0] exp__71;
  wire [9:0] wide_exponent__101;
  wire [9:0] wide_exponent__102;
  wire [9:0] exp__153;
  wire [9:0] wide_exponent__158;
  wire [9:0] wide_exponent__159;
  wire [9:0] exp__235;
  wire [9:0] wide_exponent__215;
  wire [9:0] wide_exponent__216;
  wire [9:0] exp__317;
  wire [9:0] wide_exponent__23;
  wire [7:0] high_exp__377;
  wire [22:0] result_fraction__783;
  wire [7:0] high_exp__378;
  wire [22:0] result_fraction__784;
  wire [7:0] high_exp__123;
  wire [22:0] result_fraction__522;
  wire [7:0] high_exp__124;
  wire [22:0] result_fraction__523;
  wire [9:0] wide_exponent__103;
  wire [7:0] high_exp__409;
  wire [22:0] result_fraction__816;
  wire [7:0] high_exp__410;
  wire [22:0] result_fraction__817;
  wire [7:0] high_exp__188;
  wire [22:0] result_fraction__589;
  wire [7:0] high_exp__189;
  wire [22:0] result_fraction__590;
  wire [9:0] wide_exponent__160;
  wire [7:0] high_exp__441;
  wire [22:0] result_fraction__849;
  wire [7:0] high_exp__442;
  wire [22:0] result_fraction__850;
  wire [7:0] high_exp__256;
  wire [22:0] result_fraction__656;
  wire [7:0] high_exp__257;
  wire [22:0] result_fraction__657;
  wire [9:0] wide_exponent__217;
  wire [7:0] high_exp__473;
  wire [22:0] result_fraction__882;
  wire [7:0] high_exp__474;
  wire [22:0] result_fraction__883;
  wire [7:0] high_exp__329;
  wire [22:0] result_fraction__733;
  wire [7:0] high_exp__330;
  wire [22:0] result_fraction__734;
  wire [7:0] high_exp__363;
  wire [22:0] result_fraction__768;
  wire [7:0] high_exp__364;
  wire [22:0] result_fraction__769;
  wire [7:0] high_exp__125;
  wire [22:0] result_fraction__524;
  wire [7:0] high_exp__126;
  wire [22:0] result_fraction__525;
  wire ne_169972;
  wire ne_169974;
  wire eq_169975;
  wire eq_169976;
  wire eq_169977;
  wire eq_169978;
  wire [8:0] result_exp__51;
  wire [7:0] high_exp__395;
  wire [22:0] result_fraction__801;
  wire [7:0] high_exp__396;
  wire [22:0] result_fraction__802;
  wire [7:0] high_exp__190;
  wire [22:0] result_fraction__591;
  wire [7:0] high_exp__191;
  wire [22:0] result_fraction__592;
  wire ne_169992;
  wire ne_169994;
  wire eq_169995;
  wire eq_169996;
  wire eq_169997;
  wire eq_169998;
  wire [8:0] result_exp__109;
  wire [7:0] high_exp__427;
  wire [22:0] result_fraction__834;
  wire [7:0] high_exp__428;
  wire [22:0] result_fraction__835;
  wire [7:0] high_exp__258;
  wire [22:0] result_fraction__658;
  wire [7:0] high_exp__259;
  wire [22:0] result_fraction__659;
  wire ne_170012;
  wire ne_170014;
  wire eq_170015;
  wire eq_170016;
  wire eq_170017;
  wire eq_170018;
  wire [8:0] result_exp__169;
  wire [7:0] high_exp__459;
  wire [22:0] result_fraction__867;
  wire [7:0] high_exp__460;
  wire [22:0] result_fraction__868;
  wire [7:0] high_exp__331;
  wire [22:0] result_fraction__735;
  wire [7:0] high_exp__332;
  wire [22:0] result_fraction__736;
  wire ne_170032;
  wire ne_170034;
  wire eq_170035;
  wire eq_170036;
  wire eq_170037;
  wire eq_170038;
  wire [8:0] result_exp__229;
  wire ne_170043;
  wire ne_170045;
  wire eq_170046;
  wire eq_170047;
  wire eq_170048;
  wire eq_170049;
  wire [8:0] result_exp__52;
  wire ne_170059;
  wire ne_170061;
  wire eq_170062;
  wire eq_170063;
  wire eq_170064;
  wire eq_170065;
  wire [8:0] result_exp__111;
  wire ne_170075;
  wire ne_170077;
  wire eq_170078;
  wire eq_170079;
  wire eq_170080;
  wire eq_170081;
  wire [8:0] result_exp__171;
  wire ne_170091;
  wire ne_170093;
  wire eq_170094;
  wire eq_170095;
  wire eq_170096;
  wire eq_170097;
  wire [7:0] high_exp__334;
  wire [22:0] result_fraction__738;
  wire [22:0] result_fraction__737;
  wire [8:0] result_exp__231;
  wire [8:0] wide_exponent__50;
  wire has_pos_inf__16;
  wire has_neg_inf__16;
  wire [8:0] wide_exponent__104;
  wire has_pos_inf__34;
  wire has_neg_inf__34;
  wire [8:0] wide_exponent__161;
  wire has_pos_inf__53;
  wire has_neg_inf__53;
  wire [8:0] wide_exponent__218;
  wire has_pos_inf__72;
  wire has_neg_inf__72;
  wire eq_170147;
  wire ne_170148;
  wire [8:0] wide_exponent__24;
  wire has_pos_inf__8;
  wire has_neg_inf__8;
  wire and_reduce_170162;
  wire [8:0] wide_exponent__105;
  wire has_pos_inf__35;
  wire has_neg_inf__35;
  wire and_reduce_170174;
  wire [8:0] wide_exponent__162;
  wire has_pos_inf__54;
  wire has_neg_inf__54;
  wire and_reduce_170186;
  wire [8:0] wide_exponent__219;
  wire has_pos_inf__73;
  wire has_neg_inf__73;
  wire is_result_nan__150;
  wire has_inf_arg__77;
  wire and_reduce_170200;
  wire is_result_nan__33;
  wire is_operand_inf__16;
  wire and_reduce_170214;
  wire [7:0] high_exp__129;
  wire is_result_nan__70;
  wire is_operand_inf__34;
  wire and_reduce_170230;
  wire [7:0] high_exp__194;
  wire is_result_nan__109;
  wire is_operand_inf__53;
  wire and_reduce_170246;
  wire [7:0] high_exp__262;
  wire is_result_nan__148;
  wire is_operand_inf__72;
  wire and_reduce_170262;
  wire [7:0] high_exp__336;
  wire is_result_nan__16;
  wire is_operand_inf__8;
  wire and_reduce_170270;
  wire [2:0] fraction_shift__380;
  wire [2:0] fraction_shift__255;
  wire is_subnormal__17;
  wire [7:0] high_exp__127;
  wire [7:0] result_exp__53;
  wire is_result_nan__71;
  wire is_operand_inf__35;
  wire and_reduce_170283;
  wire [2:0] fraction_shift__398;
  wire [2:0] fraction_shift__290;
  wire is_subnormal__37;
  wire [7:0] high_exp__192;
  wire [7:0] result_exp__113;
  wire is_result_nan__110;
  wire is_operand_inf__54;
  wire and_reduce_170296;
  wire [2:0] fraction_shift__416;
  wire [2:0] fraction_shift__325;
  wire is_subnormal__57;
  wire [7:0] high_exp__260;
  wire [7:0] result_exp__173;
  wire is_result_nan__149;
  wire is_operand_inf__73;
  wire and_reduce_170309;
  wire [2:0] fraction_shift__434;
  wire [2:0] fraction_shift__360;
  wire is_subnormal__77;
  wire [7:0] high_exp__333;
  wire [7:0] result_exp__233;
  wire [2:0] fraction_shift__381;
  wire [2:0] fraction_shift__256;
  wire [7:0] high_exp__128;
  wire [2:0] fraction_shift__51;
  wire result_sign__457;
  wire [7:0] result_exponent__17;
  wire result_sign__458;
  wire [2:0] fraction_shift__399;
  wire [2:0] fraction_shift__291;
  wire [7:0] high_exp__193;
  wire [2:0] fraction_shift__104;
  wire result_sign__554;
  wire [7:0] result_exponent__34;
  wire result_sign__555;
  wire [2:0] fraction_shift__417;
  wire [2:0] fraction_shift__326;
  wire [7:0] high_exp__261;
  wire [2:0] fraction_shift__161;
  wire result_sign__656;
  wire [7:0] result_exponent__53;
  wire result_sign__657;
  wire [2:0] fraction_shift__435;
  wire [2:0] fraction_shift__361;
  wire [7:0] high_exp__335;
  wire [2:0] fraction_shift__218;
  wire result_sign__768;
  wire [7:0] result_exponent__72;
  wire result_sign__769;
  wire [2:0] fraction_shift__24;
  wire result_sign__459;
  wire [7:0] result_exponent__8;
  wire [27:0] shrl_170369;
  wire [8:0] concat_170373;
  wire [2:0] fraction_shift__105;
  wire result_sign__556;
  wire [7:0] result_exponent__35;
  wire [27:0] shrl_170378;
  wire [8:0] concat_170382;
  wire [2:0] fraction_shift__162;
  wire result_sign__658;
  wire [7:0] result_exponent__54;
  wire [27:0] shrl_170387;
  wire [8:0] concat_170391;
  wire [2:0] fraction_shift__219;
  wire result_sign__770;
  wire [7:0] result_exponent__73;
  wire [27:0] shrl_170396;
  wire [8:0] concat_170400;
  wire [27:0] shrl_170401;
  wire [22:0] result_fraction__99;
  wire [22:0] result_fraction__102;
  wire [8:0] sum__17;
  wire [27:0] shrl_170409;
  wire [22:0] result_fraction__208;
  wire [22:0] result_fraction__214;
  wire [8:0] sum__36;
  wire [27:0] shrl_170417;
  wire [22:0] result_fraction__325;
  wire [22:0] result_fraction__331;
  wire [8:0] sum__55;
  wire [27:0] shrl_170425;
  wire [22:0] result_fraction__442;
  wire [22:0] result_fraction__448;
  wire [8:0] sum__74;
  wire [22:0] result_fraction__46;
  wire [8:0] sum__18;
  wire [22:0] result_fraction__100;
  wire [22:0] nan_fraction__98;
  wire [22:0] result_fraction__103;
  wire [22:0] nan_fraction__100;
  wire [22:0] result_fraction__209;
  wire [8:0] sum__37;
  wire [22:0] result_fraction__210;
  wire [22:0] nan_fraction__125;
  wire [22:0] result_fraction__216;
  wire [22:0] nan_fraction__127;
  wire [22:0] result_fraction__326;
  wire [8:0] sum__56;
  wire [22:0] result_fraction__327;
  wire [22:0] nan_fraction__154;
  wire [22:0] result_fraction__333;
  wire [22:0] nan_fraction__156;
  wire [22:0] result_fraction__443;
  wire [8:0] sum__75;
  wire [22:0] result_fraction__444;
  wire [22:0] nan_fraction__183;
  wire [22:0] result_fraction__450;
  wire [22:0] nan_fraction__185;
  wire [22:0] result_fraction__47;
  wire [22:0] nan_fraction__99;
  wire [22:0] result_fraction__101;
  wire [22:0] result_fraction__104;
  wire [7:0] prod_bexp__70;
  wire [7:0] x_bexp__796;
  wire [22:0] result_fraction__211;
  wire [22:0] nan_fraction__126;
  wire [22:0] result_fraction__212;
  wire [22:0] result_fraction__218;
  wire [7:0] prod_bexp__139;
  wire [7:0] x_bexp__797;
  wire [22:0] result_fraction__328;
  wire [22:0] nan_fraction__155;
  wire [22:0] result_fraction__329;
  wire [22:0] result_fraction__335;
  wire [7:0] prod_bexp__211;
  wire [7:0] x_bexp__798;
  wire [22:0] result_fraction__445;
  wire [22:0] nan_fraction__184;
  wire [22:0] result_fraction__446;
  wire [22:0] result_fraction__452;
  wire [7:0] prod_bexp__283;
  wire [7:0] x_bexp__799;
  wire [22:0] result_fraction__48;
  wire [7:0] prod_bexp__34;
  wire [7:0] x_bexp__800;
  wire fraction_is_zero__16;
  wire [22:0] prod_fraction__51;
  wire [7:0] incremented_sum__92;
  wire [22:0] result_fraction__213;
  wire [7:0] prod_bexp__140;
  wire [7:0] x_bexp__801;
  wire fraction_is_zero__34;
  wire [22:0] prod_fraction__103;
  wire [7:0] incremented_sum__110;
  wire [22:0] result_fraction__330;
  wire [7:0] prod_bexp__212;
  wire [7:0] x_bexp__802;
  wire fraction_is_zero__53;
  wire [22:0] prod_fraction__157;
  wire [7:0] incremented_sum__128;
  wire [22:0] result_fraction__447;
  wire [7:0] prod_bexp__284;
  wire [7:0] x_bexp__803;
  wire fraction_is_zero__72;
  wire [22:0] prod_fraction__211;
  wire [7:0] incremented_sum__146;
  wire fraction_is_zero__8;
  wire [22:0] prod_fraction__25;
  wire [7:0] incremented_sum__93;
  wire [27:0] wide_y__34;
  wire [7:0] x_bexpbs_difference__18;
  wire fraction_is_zero__35;
  wire [22:0] prod_fraction__104;
  wire [7:0] incremented_sum__111;
  wire [27:0] wide_y__71;
  wire [7:0] x_bexpbs_difference__35;
  wire fraction_is_zero__54;
  wire [22:0] prod_fraction__158;
  wire [7:0] incremented_sum__129;
  wire [27:0] wide_y__109;
  wire [7:0] x_bexpbs_difference__53;
  wire fraction_is_zero__73;
  wire [22:0] prod_fraction__212;
  wire [7:0] incremented_sum__147;
  wire [27:0] wide_y__147;
  wire [7:0] x_bexpbs_difference__71;
  wire [27:0] wide_y__17;
  wire [7:0] x_bexpbs_difference__9;
  wire [2:0] concat_170634;
  wire [7:0] x_bexp__142;
  wire [7:0] x_bexp__804;
  wire [27:0] wide_y__35;
  wire [7:0] sub_170640;
  wire [27:0] wide_y__72;
  wire [7:0] x_bexpbs_difference__36;
  wire [2:0] concat_170646;
  wire [7:0] x_bexp__283;
  wire [7:0] x_bexp__805;
  wire [27:0] wide_y__73;
  wire [7:0] sub_170652;
  wire [27:0] wide_y__110;
  wire [7:0] x_bexpbs_difference__54;
  wire [2:0] concat_170658;
  wire [7:0] x_bexp__427;
  wire [7:0] x_bexp__806;
  wire [27:0] wide_y__111;
  wire [7:0] sub_170664;
  wire [27:0] wide_y__148;
  wire [7:0] x_bexpbs_difference__72;
  wire [2:0] concat_170670;
  wire [7:0] x_bexp__571;
  wire [7:0] x_bexp__807;
  wire [27:0] wide_y__149;
  wire [7:0] sub_170676;
  wire [2:0] concat_170677;
  wire [7:0] x_bexp__70;
  wire [7:0] x_bexp__808;
  wire [27:0] wide_y__36;
  wire [7:0] sub_170683;
  wire result_sign__82;
  wire [22:0] x_fraction__142;
  wire [27:0] dropped__17;
  wire [2:0] concat_170691;
  wire [7:0] x_bexp__284;
  wire [7:0] x_bexp__809;
  wire [27:0] wide_y__74;
  wire [7:0] sub_170697;
  wire result_sign__172;
  wire [22:0] x_fraction__283;
  wire [27:0] dropped__36;
  wire [2:0] concat_170705;
  wire [7:0] x_bexp__428;
  wire [7:0] x_bexp__810;
  wire [27:0] wide_y__112;
  wire [7:0] sub_170711;
  wire result_sign__269;
  wire [22:0] x_fraction__427;
  wire [27:0] dropped__55;
  wire [2:0] concat_170719;
  wire [7:0] x_bexp__572;
  wire [7:0] x_bexp__811;
  wire [27:0] wide_y__150;
  wire [7:0] sub_170725;
  wire result_sign__366;
  wire [22:0] x_fraction__571;
  wire [27:0] dropped__74;
  wire result_sign__38;
  wire [22:0] x_fraction__70;
  wire [27:0] dropped__18;
  wire result_sign__83;
  wire [27:0] wide_x__34;
  wire result_sign__173;
  wire [22:0] x_fraction__284;
  wire [27:0] dropped__37;
  wire result_sign__174;
  wire [27:0] wide_x__71;
  wire result_sign__270;
  wire [22:0] x_fraction__428;
  wire [27:0] dropped__56;
  wire result_sign__271;
  wire [27:0] wide_x__109;
  wire result_sign__367;
  wire [22:0] x_fraction__572;
  wire [27:0] dropped__75;
  wire x_sign__141;
  wire result_sign__368;
  wire [27:0] wide_x__147;
  wire result_sign__39;
  wire [27:0] wide_x__17;
  wire result_sign__84;
  wire [27:0] wide_x__35;
  wire result_sign__175;
  wire [27:0] wide_x__72;
  wire result_sign__176;
  wire [27:0] wide_x__73;
  wire result_sign__272;
  wire [27:0] wide_x__110;
  wire result_sign__273;
  wire [27:0] wide_x__111;
  wire result_sign__369;
  wire [27:0] wide_x__148;
  wire result_sign__374;
  wire result_sign__370;
  wire [27:0] wide_x__149;
  wire result_sign__40;
  wire [27:0] wide_x__36;
  wire x_sign__36;
  wire prod_sign__17;
  wire [27:0] neg_170834;
  wire [27:0] sticky__53;
  wire result_sign__177;
  wire [27:0] wide_x__74;
  wire x_sign__71;
  wire prod_sign__35;
  wire [27:0] neg_170843;
  wire [27:0] sticky__112;
  wire result_sign__274;
  wire [27:0] wide_x__112;
  wire x_sign__107;
  wire prod_sign__53;
  wire [27:0] neg_170852;
  wire [27:0] sticky__171;
  wire result_sign__371;
  wire [27:0] wide_x__150;
  wire x_sign__143;
  wire prod_sign__71;
  wire [27:0] neg_170861;
  wire [27:0] sticky__230;
  wire x_sign__18;
  wire prod_sign__18;
  wire [27:0] neg_170866;
  wire [27:0] sticky__54;
  wire [27:0] xddend_y__17;
  wire x_sign__72;
  wire prod_sign__36;
  wire [27:0] neg_170875;
  wire [27:0] sticky__113;
  wire [27:0] xddend_y__35;
  wire x_sign__108;
  wire prod_sign__54;
  wire [27:0] neg_170884;
  wire [27:0] sticky__172;
  wire [27:0] xddend_y__53;
  wire x_sign__144;
  wire prod_sign__72;
  wire [27:0] neg_170893;
  wire [27:0] sticky__231;
  wire [27:0] xddend_y__71;
  wire [27:0] xddend_y__18;
  wire [24:0] sel_170904;
  wire result_sign__1084;
  wire [27:0] xddend_y__36;
  wire [24:0] sel_170911;
  wire result_sign__1085;
  wire [27:0] xddend_y__54;
  wire [24:0] sel_170918;
  wire result_sign__1086;
  wire [27:0] xddend_y__72;
  wire [24:0] sel_170925;
  wire result_sign__1087;
  wire [24:0] sel_170928;
  wire result_sign__1088;
  wire [24:0] sel_170933;
  wire result_sign__1089;
  wire [24:0] sel_170938;
  wire result_sign__1090;
  wire [24:0] sel_170943;
  wire result_sign__1091;
  wire [25:0] add_170950;
  wire [25:0] add_170953;
  wire [25:0] add_170956;
  wire [25:0] add_170959;
  wire [25:0] add_170960;
  wire [25:0] add_170963;
  wire [25:0] add_170966;
  wire [25:0] add_170969;
  wire [27:0] concat_170974;
  wire [27:0] concat_170977;
  wire [27:0] concat_170980;
  wire [27:0] concat_170983;
  wire [27:0] concat_170984;
  wire [27:0] concat_170987;
  wire [27:0] concat_170990;
  wire [27:0] concat_170993;
  wire [27:0] xbs_fraction__17;
  wire [27:0] xbs_fraction__35;
  wire [27:0] xbs_fraction__53;
  wire [27:0] xbs_fraction__71;
  wire [27:0] xbs_fraction__18;
  wire [27:0] reverse_171009;
  wire [27:0] xbs_fraction__36;
  wire [27:0] reverse_171011;
  wire [27:0] xbs_fraction__54;
  wire [27:0] reverse_171013;
  wire [27:0] xbs_fraction__72;
  wire [27:0] reverse_171015;
  wire [27:0] reverse_171016;
  wire [28:0] one_hot_171017;
  wire [27:0] reverse_171018;
  wire [28:0] one_hot_171019;
  wire [27:0] reverse_171020;
  wire [28:0] one_hot_171021;
  wire [27:0] reverse_171022;
  wire [28:0] one_hot_171023;
  wire [28:0] one_hot_171024;
  wire [4:0] encode_171025;
  wire [28:0] one_hot_171026;
  wire [4:0] encode_171027;
  wire [28:0] one_hot_171028;
  wire [4:0] encode_171029;
  wire [28:0] one_hot_171030;
  wire [4:0] encode_171031;
  wire [4:0] encode_171032;
  wire [4:0] encode_171034;
  wire [4:0] encode_171036;
  wire [4:0] encode_171038;
  wire cancel__18;
  wire carry_bit__17;
  wire [22:0] result_fraction__526;
  wire cancel__36;
  wire carry_bit__36;
  wire [22:0] result_fraction__593;
  wire cancel__55;
  wire carry_bit__55;
  wire [22:0] result_fraction__660;
  wire cancel__74;
  wire carry_bit__74;
  wire [22:0] result_fraction__739;
  wire cancel__9;
  wire carry_bit__18;
  wire [22:0] result_fraction__527;
  wire [27:0] leading_zeroes__17;
  wire cancel__37;
  wire carry_bit__37;
  wire [22:0] result_fraction__594;
  wire [27:0] leading_zeroes__36;
  wire cancel__56;
  wire carry_bit__56;
  wire [22:0] result_fraction__661;
  wire [27:0] leading_zeroes__55;
  wire cancel__75;
  wire carry_bit__75;
  wire [22:0] result_fraction__740;
  wire [27:0] leading_zeroes__74;
  wire [27:0] leading_zeroes__18;
  wire [26:0] carry_fraction__34;
  wire [27:0] add_171104;
  wire [27:0] leading_zeroes__37;
  wire [26:0] carry_fraction__71;
  wire [27:0] add_171117;
  wire [27:0] leading_zeroes__56;
  wire [26:0] carry_fraction__109;
  wire [27:0] add_171130;
  wire [27:0] leading_zeroes__75;
  wire [26:0] carry_fraction__147;
  wire [27:0] add_171143;
  wire [26:0] carry_fraction__17;
  wire [27:0] add_171150;
  wire [2:0] concat_171151;
  wire [26:0] carry_fraction__35;
  wire [26:0] cancel_fraction__17;
  wire [26:0] carry_fraction__72;
  wire [27:0] add_171160;
  wire [2:0] concat_171161;
  wire [26:0] carry_fraction__73;
  wire [26:0] cancel_fraction__36;
  wire [26:0] carry_fraction__110;
  wire [27:0] add_171170;
  wire [2:0] concat_171171;
  wire [26:0] carry_fraction__111;
  wire [26:0] cancel_fraction__55;
  wire [26:0] carry_fraction__148;
  wire [27:0] add_171180;
  wire [2:0] concat_171181;
  wire [26:0] carry_fraction__149;
  wire [26:0] cancel_fraction__74;
  wire [2:0] concat_171184;
  wire [26:0] carry_fraction__36;
  wire [26:0] cancel_fraction__18;
  wire [26:0] shifted_fraction__17;
  wire [2:0] concat_171188;
  wire [26:0] carry_fraction__74;
  wire [26:0] cancel_fraction__37;
  wire [26:0] shifted_fraction__36;
  wire [2:0] concat_171192;
  wire [26:0] carry_fraction__112;
  wire [26:0] cancel_fraction__56;
  wire [26:0] shifted_fraction__55;
  wire [2:0] concat_171196;
  wire [26:0] carry_fraction__150;
  wire [26:0] cancel_fraction__75;
  wire [26:0] shifted_fraction__74;
  wire [26:0] shifted_fraction__18;
  wire result_sign__1092;
  wire [26:0] shifted_fraction__37;
  wire result_sign__1093;
  wire [26:0] shifted_fraction__56;
  wire result_sign__1094;
  wire [26:0] shifted_fraction__75;
  wire result_sign__1095;
  wire result_sign__1096;
  wire [2:0] normal_chunk__17;
  wire [2:0] fraction_shift__257;
  wire [1:0] half_way_chunk__17;
  wire result_sign__1097;
  wire [2:0] normal_chunk__36;
  wire [2:0] fraction_shift__292;
  wire [1:0] half_way_chunk__36;
  wire result_sign__1098;
  wire [2:0] normal_chunk__55;
  wire [2:0] fraction_shift__327;
  wire [1:0] half_way_chunk__55;
  wire result_sign__1099;
  wire [2:0] normal_chunk__74;
  wire [2:0] fraction_shift__362;
  wire [1:0] half_way_chunk__74;
  wire [2:0] normal_chunk__18;
  wire [2:0] fraction_shift__258;
  wire [1:0] half_way_chunk__18;
  wire result_sign__460;
  wire [24:0] add_171253;
  wire [2:0] normal_chunk__37;
  wire [2:0] fraction_shift__293;
  wire [1:0] half_way_chunk__37;
  wire result_sign__557;
  wire [24:0] add_171263;
  wire [2:0] normal_chunk__56;
  wire [2:0] fraction_shift__328;
  wire [1:0] half_way_chunk__56;
  wire result_sign__659;
  wire [24:0] add_171273;
  wire [2:0] normal_chunk__75;
  wire [2:0] fraction_shift__363;
  wire [1:0] half_way_chunk__75;
  wire result_sign__771;
  wire [24:0] add_171283;
  wire result_sign__461;
  wire [24:0] add_171287;
  wire do_round_up__35;
  wire result_sign__558;
  wire [24:0] add_171294;
  wire do_round_up__74;
  wire result_sign__660;
  wire [24:0] add_171301;
  wire do_round_up__113;
  wire result_sign__772;
  wire [24:0] add_171308;
  wire do_round_up__152;
  wire do_round_up__36;
  wire [27:0] rounded_fraction__17;
  wire do_round_up__75;
  wire [27:0] rounded_fraction__36;
  wire do_round_up__114;
  wire [27:0] rounded_fraction__55;
  wire do_round_up__153;
  wire [27:0] rounded_fraction__74;
  wire [27:0] rounded_fraction__18;
  wire result_sign__462;
  wire [7:0] x_bexp__590;
  wire rounding_carry__17;
  wire [27:0] rounded_fraction__37;
  wire result_sign__559;
  wire [7:0] x_bexp__608;
  wire rounding_carry__36;
  wire [27:0] rounded_fraction__56;
  wire result_sign__661;
  wire [7:0] x_bexp__626;
  wire rounding_carry__55;
  wire [27:0] rounded_fraction__75;
  wire result_sign__773;
  wire [7:0] x_bexp__644;
  wire rounding_carry__74;
  wire result_sign__463;
  wire [7:0] x_bexp__591;
  wire rounding_carry__18;
  wire result_sign__560;
  wire [7:0] x_bexp__609;
  wire rounding_carry__37;
  wire result_sign__662;
  wire [7:0] x_bexp__627;
  wire rounding_carry__56;
  wire result_sign__774;
  wire [7:0] x_bexp__645;
  wire rounding_carry__75;
  wire result_sign__464;
  wire [8:0] add_171367;
  wire result_sign__561;
  wire [8:0] add_171373;
  wire result_sign__663;
  wire [8:0] add_171379;
  wire result_sign__775;
  wire [8:0] add_171385;
  wire result_sign__465;
  wire [8:0] add_171389;
  wire result_sign__562;
  wire [8:0] add_171398;
  wire result_sign__664;
  wire [8:0] add_171407;
  wire result_sign__776;
  wire [8:0] add_171416;
  wire [9:0] add_171429;
  wire [9:0] add_171437;
  wire [9:0] add_171445;
  wire [9:0] add_171453;
  wire [9:0] add_171456;
  wire [9:0] wide_exponent__51;
  wire [9:0] add_171461;
  wire [9:0] wide_exponent__106;
  wire [9:0] add_171466;
  wire [9:0] wide_exponent__163;
  wire [9:0] add_171471;
  wire [9:0] wide_exponent__220;
  wire [9:0] wide_exponent__25;
  wire [9:0] wide_exponent__52;
  wire [9:0] wide_exponent__107;
  wire [9:0] wide_exponent__108;
  wire [9:0] wide_exponent__164;
  wire [9:0] wide_exponent__165;
  wire [9:0] wide_exponent__221;
  wire [9:0] wide_exponent__222;
  wire [9:0] wide_exponent__26;
  wire [9:0] wide_exponent__109;
  wire [9:0] wide_exponent__166;
  wire [9:0] wide_exponent__223;
  wire [7:0] high_exp__130;
  wire [22:0] result_fraction__528;
  wire [7:0] high_exp__131;
  wire [22:0] result_fraction__529;
  wire [8:0] wide_exponent__53;
  wire [7:0] high_exp__195;
  wire [22:0] result_fraction__595;
  wire [7:0] high_exp__196;
  wire [22:0] result_fraction__596;
  wire [8:0] wide_exponent__110;
  wire [7:0] high_exp__263;
  wire [22:0] result_fraction__662;
  wire [7:0] high_exp__264;
  wire [22:0] result_fraction__663;
  wire [8:0] wide_exponent__167;
  wire [7:0] high_exp__337;
  wire [22:0] result_fraction__741;
  wire [7:0] high_exp__338;
  wire [22:0] result_fraction__742;
  wire [8:0] wide_exponent__224;
  wire [7:0] high_exp__132;
  wire [22:0] result_fraction__530;
  wire [7:0] high_exp__133;
  wire [22:0] result_fraction__531;
  wire [8:0] wide_exponent__54;
  wire eq_171549;
  wire eq_171550;
  wire eq_171551;
  wire eq_171552;
  wire [7:0] high_exp__381;
  wire [22:0] result_fraction__787;
  wire [7:0] high_exp__382;
  wire [22:0] result_fraction__788;
  wire [7:0] high_exp__197;
  wire [22:0] result_fraction__597;
  wire [7:0] high_exp__198;
  wire [22:0] result_fraction__598;
  wire [8:0] wide_exponent__111;
  wire eq_171563;
  wire eq_171564;
  wire eq_171565;
  wire eq_171566;
  wire [7:0] high_exp__413;
  wire [22:0] result_fraction__820;
  wire [7:0] high_exp__414;
  wire [22:0] result_fraction__821;
  wire [7:0] high_exp__265;
  wire [22:0] result_fraction__664;
  wire [7:0] high_exp__266;
  wire [22:0] result_fraction__665;
  wire [8:0] wide_exponent__168;
  wire eq_171577;
  wire eq_171578;
  wire eq_171579;
  wire eq_171580;
  wire [7:0] high_exp__445;
  wire [22:0] result_fraction__853;
  wire [7:0] high_exp__446;
  wire [22:0] result_fraction__854;
  wire [7:0] high_exp__339;
  wire [22:0] result_fraction__743;
  wire [7:0] high_exp__340;
  wire [22:0] result_fraction__744;
  wire [8:0] wide_exponent__225;
  wire eq_171591;
  wire eq_171592;
  wire eq_171593;
  wire eq_171594;
  wire [7:0] high_exp__477;
  wire [22:0] result_fraction__886;
  wire [7:0] high_exp__478;
  wire [22:0] result_fraction__887;
  wire eq_171600;
  wire eq_171601;
  wire eq_171602;
  wire eq_171603;
  wire [7:0] high_exp__379;
  wire [22:0] result_fraction__785;
  wire [7:0] high_exp__380;
  wire [22:0] result_fraction__786;
  wire ne_171615;
  wire ne_171617;
  wire eq_171618;
  wire eq_171619;
  wire eq_171620;
  wire eq_171621;
  wire [7:0] high_exp__411;
  wire [22:0] result_fraction__818;
  wire [7:0] high_exp__412;
  wire [22:0] result_fraction__819;
  wire ne_171633;
  wire ne_171635;
  wire eq_171636;
  wire eq_171637;
  wire eq_171638;
  wire eq_171639;
  wire [7:0] high_exp__443;
  wire [22:0] result_fraction__851;
  wire [7:0] high_exp__444;
  wire [22:0] result_fraction__852;
  wire ne_171651;
  wire ne_171653;
  wire eq_171654;
  wire eq_171655;
  wire eq_171656;
  wire eq_171657;
  wire [7:0] high_exp__475;
  wire [22:0] result_fraction__884;
  wire [7:0] high_exp__476;
  wire [22:0] result_fraction__885;
  wire ne_171669;
  wire ne_171671;
  wire ne_171678;
  wire ne_171680;
  wire [2:0] fraction_shift__382;
  wire [2:0] fraction_shift__259;
  wire is_operand_inf__17;
  wire and_reduce_171685;
  wire ne_171697;
  wire ne_171699;
  wire [2:0] fraction_shift__400;
  wire [2:0] fraction_shift__294;
  wire is_operand_inf__36;
  wire and_reduce_171704;
  wire ne_171716;
  wire ne_171718;
  wire [2:0] fraction_shift__418;
  wire [2:0] fraction_shift__329;
  wire is_operand_inf__55;
  wire and_reduce_171723;
  wire ne_171735;
  wire ne_171737;
  wire [2:0] fraction_shift__436;
  wire [2:0] fraction_shift__364;
  wire is_operand_inf__74;
  wire and_reduce_171742;
  wire [2:0] fraction_shift__383;
  wire [2:0] fraction_shift__260;
  wire is_operand_inf__18;
  wire and_reduce_171752;
  wire [2:0] fraction_shift__54;
  wire has_pos_inf__17;
  wire has_neg_inf__17;
  wire [2:0] fraction_shift__401;
  wire [2:0] fraction_shift__295;
  wire is_operand_inf__37;
  wire and_reduce_171766;
  wire [2:0] fraction_shift__110;
  wire has_pos_inf__36;
  wire has_neg_inf__36;
  wire [2:0] fraction_shift__419;
  wire [2:0] fraction_shift__330;
  wire is_operand_inf__56;
  wire and_reduce_171780;
  wire [2:0] fraction_shift__167;
  wire has_pos_inf__55;
  wire has_neg_inf__55;
  wire [2:0] fraction_shift__437;
  wire [2:0] fraction_shift__365;
  wire is_operand_inf__75;
  wire and_reduce_171794;
  wire [2:0] fraction_shift__224;
  wire has_pos_inf__74;
  wire has_neg_inf__74;
  wire [2:0] fraction_shift__27;
  wire has_pos_inf__18;
  wire has_neg_inf__18;
  wire [27:0] shrl_171808;
  wire [2:0] fraction_shift__111;
  wire has_pos_inf__37;
  wire has_neg_inf__37;
  wire [27:0] shrl_171817;
  wire [2:0] fraction_shift__168;
  wire has_pos_inf__56;
  wire has_neg_inf__56;
  wire [27:0] shrl_171826;
  wire [2:0] fraction_shift__225;
  wire has_pos_inf__75;
  wire has_neg_inf__75;
  wire [27:0] shrl_171835;
  wire [27:0] shrl_171840;
  wire [22:0] result_fraction__105;
  wire is_result_nan__35;
  wire [27:0] shrl_171848;
  wire [22:0] result_fraction__220;
  wire is_result_nan__74;
  wire [27:0] shrl_171856;
  wire [22:0] result_fraction__337;
  wire is_result_nan__113;
  wire [27:0] shrl_171864;
  wire [22:0] result_fraction__454;
  wire is_result_nan__152;
  wire [22:0] result_fraction__52;
  wire is_result_nan__36;
  wire [22:0] result_fraction__106;
  wire [22:0] nan_fraction__101;
  wire or_171877;
  wire [7:0] high_exp__134;
  wire [22:0] result_fraction__221;
  wire is_result_nan__75;
  wire [22:0] result_fraction__222;
  wire [22:0] nan_fraction__128;
  wire [7:0] high_exp__199;
  wire [22:0] result_fraction__338;
  wire is_result_nan__114;
  wire [22:0] result_fraction__339;
  wire [22:0] nan_fraction__157;
  wire [7:0] high_exp__267;
  wire [22:0] result_fraction__455;
  wire is_result_nan__153;
  wire [22:0] result_fraction__456;
  wire [22:0] nan_fraction__186;
  wire [7:0] high_exp__341;
  wire [22:0] result_fraction__53;
  wire [22:0] nan_fraction__102;
  wire or_171902;
  wire [7:0] high_exp__135;
  wire result_sign__466;
  wire [22:0] result_fraction__107;
  wire [7:0] result_exponent__18;
  wire [7:0] x_bexp__812;
  wire [22:0] result_fraction__223;
  wire [22:0] nan_fraction__129;
  wire or_171910;
  wire [7:0] high_exp__200;
  wire result_sign__563;
  wire [22:0] result_fraction__224;
  wire [7:0] result_exponent__36;
  wire [7:0] x_bexp__813;
  wire [22:0] result_fraction__340;
  wire [22:0] nan_fraction__158;
  wire or_171918;
  wire [7:0] high_exp__268;
  wire result_sign__665;
  wire [22:0] result_fraction__341;
  wire [7:0] result_exponent__55;
  wire [7:0] x_bexp__814;
  wire [22:0] result_fraction__457;
  wire [22:0] nan_fraction__187;
  wire or_171926;
  wire [7:0] high_exp__342;
  wire result_sign__777;
  wire [22:0] result_fraction__458;
  wire [7:0] result_exponent__74;
  wire [7:0] x_bexp__815;
  wire result_sign__467;
  wire [22:0] result_fraction__108;
  wire [7:0] result_exponent__9;
  wire [7:0] x_bexp__816;
  wire ne_171938;
  wire result_sign__564;
  wire [22:0] result_fraction__225;
  wire [7:0] result_exponent__37;
  wire [7:0] x_bexp__817;
  wire ne_171945;
  wire result_sign__666;
  wire [22:0] result_fraction__342;
  wire [7:0] result_exponent__56;
  wire [7:0] x_bexp__818;
  wire ne_171952;
  wire result_sign__778;
  wire [22:0] result_fraction__459;
  wire [7:0] result_exponent__75;
  wire [7:0] x_bexp__819;
  wire ne_171959;
  wire ne_171962;
  wire result_sign__468;
  wire [23:0] y_stencil_out_fraction__5;
  wire ne_171968;
  wire result_sign__565;
  wire [23:0] y_stencil_out_fraction__13;
  wire ne_171974;
  wire result_sign__667;
  wire [23:0] y_stencil_out_fraction__23;
  wire ne_171980;
  wire result_sign__779;
  wire [23:0] y_stencil_out_fraction__33;
  wire result_sign__469;
  wire [23:0] x_stencil_out_fraction__5;
  wire [23:0] y_stencil_out_fraction__3;
  wire result_sign__566;
  wire [23:0] x_stencil_out_fraction__13;
  wire [23:0] y_stencil_out_fraction__15;
  wire result_sign__668;
  wire [23:0] x_stencil_out_fraction__23;
  wire [23:0] y_stencil_out_fraction__25;
  wire result_sign__780;
  wire [23:0] x_stencil_out_fraction__33;
  wire [23:0] y_stencil_out_fraction__35;
  wire [23:0] x_stencil_out_fraction__3;
  wire result_sign__470;
  wire [8:0] add_172007;
  wire [47:0] fraction__170;
  wire [23:0] x_stencil_out_fraction__15;
  wire result_sign__567;
  wire [8:0] add_172012;
  wire [47:0] fraction__342;
  wire [23:0] x_stencil_out_fraction__25;
  wire result_sign__669;
  wire [8:0] add_172017;
  wire [47:0] fraction__521;
  wire [23:0] x_stencil_out_fraction__35;
  wire result_sign__781;
  wire [8:0] add_172022;
  wire [47:0] fraction__700;
  wire result_sign__471;
  wire [8:0] add_172025;
  wire [47:0] fraction__163;
  wire result_sign__568;
  wire [8:0] add_172033;
  wire [47:0] fraction__343;
  wire result_sign__670;
  wire [8:0] add_172041;
  wire [47:0] fraction__522;
  wire result_sign__782;
  wire [8:0] add_172049;
  wire [47:0] fraction__701;
  wire [9:0] exp__76;
  wire [47:0] fraction__171;
  wire [47:0] sticky__56;
  wire [9:0] exp__155;
  wire [47:0] fraction__344;
  wire [47:0] sticky__114;
  wire [9:0] exp__237;
  wire [47:0] fraction__523;
  wire [47:0] sticky__173;
  wire [9:0] exp__319;
  wire [47:0] fraction__702;
  wire [47:0] sticky__232;
  wire [9:0] exp__73;
  wire [47:0] fraction__164;
  wire [47:0] sticky__55;
  wire [9:0] exp__77;
  wire [47:0] fraction__172;
  wire [9:0] exp__156;
  wire [47:0] fraction__345;
  wire [47:0] sticky__115;
  wire [9:0] exp__157;
  wire [47:0] fraction__346;
  wire [9:0] exp__238;
  wire [47:0] fraction__524;
  wire [47:0] sticky__174;
  wire [9:0] exp__239;
  wire [47:0] fraction__525;
  wire [9:0] exp__320;
  wire [47:0] fraction__703;
  wire [47:0] sticky__233;
  wire [9:0] exp__321;
  wire [47:0] fraction__704;
  wire [9:0] exp__74;
  wire [47:0] fraction__165;
  wire [9:0] exp__78;
  wire result_sign__472;
  wire [9:0] exp__158;
  wire [47:0] fraction__347;
  wire [9:0] exp__159;
  wire result_sign__569;
  wire [9:0] exp__240;
  wire [47:0] fraction__526;
  wire [9:0] exp__241;
  wire result_sign__671;
  wire [9:0] exp__322;
  wire [47:0] fraction__705;
  wire [9:0] exp__323;
  wire result_sign__783;
  wire [9:0] exp__75;
  wire result_sign__473;
  wire [9:0] exp__160;
  wire result_sign__570;
  wire [9:0] exp__242;
  wire result_sign__672;
  wire [9:0] exp__324;
  wire result_sign__784;
  wire [47:0] fraction__173;
  wire [47:0] sticky__57;
  wire [47:0] fraction__348;
  wire [47:0] sticky__116;
  wire [47:0] fraction__527;
  wire [47:0] sticky__175;
  wire [47:0] fraction__706;
  wire [47:0] sticky__234;
  wire [47:0] fraction__166;
  wire [47:0] sticky__58;
  wire [47:0] fraction__174;
  wire [47:0] fraction__349;
  wire [47:0] sticky__117;
  wire [47:0] fraction__350;
  wire [47:0] fraction__528;
  wire [47:0] sticky__176;
  wire [47:0] fraction__529;
  wire [47:0] fraction__707;
  wire [47:0] sticky__235;
  wire [47:0] fraction__708;
  wire [47:0] fraction__167;
  wire [47:0] fraction__351;
  wire [47:0] fraction__530;
  wire [47:0] fraction__709;
  wire result_sign__474;
  wire [22:0] fraction__175;
  wire result_sign__571;
  wire [22:0] fraction__352;
  wire result_sign__673;
  wire [22:0] fraction__531;
  wire result_sign__785;
  wire [22:0] fraction__710;
  wire result_sign__475;
  wire [22:0] fraction__168;
  wire greater_than_half_way__19;
  wire [23:0] fraction__176;
  wire result_sign__572;
  wire [22:0] fraction__353;
  wire greater_than_half_way__39;
  wire [23:0] fraction__354;
  wire result_sign__674;
  wire [22:0] fraction__532;
  wire greater_than_half_way__59;
  wire [23:0] fraction__533;
  wire result_sign__786;
  wire [22:0] fraction__711;
  wire greater_than_half_way__79;
  wire [23:0] fraction__712;
  wire greater_than_half_way__20;
  wire [23:0] fraction__169;
  wire do_round_up__37;
  wire [23:0] add_172321;
  wire greater_than_half_way__40;
  wire [23:0] fraction__355;
  wire do_round_up__76;
  wire [23:0] add_172327;
  wire greater_than_half_way__60;
  wire [23:0] fraction__534;
  wire do_round_up__115;
  wire [23:0] add_172333;
  wire greater_than_half_way__80;
  wire [23:0] fraction__713;
  wire do_round_up__154;
  wire [23:0] add_172339;
  wire do_round_up__38;
  wire [23:0] add_172341;
  wire [23:0] fraction__177;
  wire do_round_up__77;
  wire [23:0] add_172345;
  wire [23:0] fraction__356;
  wire do_round_up__116;
  wire [23:0] add_172349;
  wire [23:0] fraction__535;
  wire do_round_up__155;
  wire [23:0] add_172353;
  wire [23:0] fraction__714;
  wire [23:0] fraction__178;
  wire [9:0] add_172359;
  wire [23:0] fraction__357;
  wire [9:0] add_172363;
  wire [23:0] fraction__536;
  wire [9:0] add_172367;
  wire [23:0] fraction__715;
  wire [9:0] add_172371;
  wire [9:0] add_172373;
  wire [9:0] exp__79;
  wire [9:0] add_172377;
  wire [9:0] exp__161;
  wire [9:0] add_172381;
  wire [9:0] exp__243;
  wire [9:0] add_172385;
  wire [9:0] exp__325;
  wire [9:0] exp__80;
  wire [9:0] exp__162;
  wire [9:0] exp__244;
  wire [9:0] exp__326;
  wire [8:0] result_exp__57;
  wire [8:0] result_exp__115;
  wire [8:0] result_exp__175;
  wire [8:0] result_exp__235;
  wire [8:0] result_exp__55;
  wire [22:0] result_fraction__534;
  wire [22:0] result_fraction__532;
  wire [8:0] result_exp__58;
  wire [8:0] result_exp__116;
  wire [7:0] high_exp__201;
  wire [22:0] result_fraction__601;
  wire [22:0] result_fraction__599;
  wire [8:0] result_exp__117;
  wire [8:0] result_exp__176;
  wire [7:0] high_exp__269;
  wire [22:0] result_fraction__668;
  wire [22:0] result_fraction__666;
  wire [8:0] result_exp__177;
  wire [8:0] result_exp__236;
  wire [7:0] high_exp__343;
  wire [22:0] result_fraction__747;
  wire [22:0] result_fraction__745;
  wire [8:0] result_exp__237;
  wire [22:0] result_fraction__535;
  wire [22:0] result_fraction__533;
  wire [8:0] result_exp__56;
  wire [22:0] result_fraction__602;
  wire [22:0] result_fraction__600;
  wire [8:0] result_exp__118;
  wire eq_172444;
  wire [22:0] result_fraction__669;
  wire [22:0] result_fraction__667;
  wire [8:0] result_exp__178;
  wire eq_172451;
  wire [22:0] result_fraction__748;
  wire [22:0] result_fraction__746;
  wire [8:0] result_exp__238;
  wire eq_172458;
  wire is_result_nan__37;
  wire has_inf_arg__19;
  wire and_reduce_172468;
  wire is_result_nan__76;
  wire has_inf_arg__39;
  wire and_reduce_172475;
  wire is_result_nan__115;
  wire has_inf_arg__59;
  wire and_reduce_172482;
  wire is_result_nan__154;
  wire has_inf_arg__79;
  wire and_reduce_172489;
  wire is_result_nan__38;
  wire has_inf_arg__20;
  wire and_reduce_172495;
  wire [7:0] high_exp__136;
  wire is_result_nan__77;
  wire has_inf_arg__40;
  wire and_reduce_172503;
  wire [7:0] high_exp__202;
  wire is_result_nan__116;
  wire has_inf_arg__60;
  wire and_reduce_172511;
  wire [7:0] high_exp__270;
  wire is_result_nan__155;
  wire has_inf_arg__80;
  wire and_reduce_172519;
  wire [7:0] high_exp__344;
  wire is_subnormal__20;
  wire is_subnormal__19;
  wire [7:0] high_exp__137;
  wire [7:0] result_exp__59;
  wire is_subnormal__40;
  wire is_subnormal__39;
  wire [7:0] high_exp__203;
  wire [7:0] result_exp__119;
  wire is_subnormal__60;
  wire is_subnormal__59;
  wire [7:0] high_exp__271;
  wire [7:0] result_exp__179;
  wire is_subnormal__80;
  wire is_subnormal__79;
  wire [7:0] high_exp__345;
  wire [7:0] result_exp__239;
  wire result_sign__476;
  wire [7:0] result_exp__60;
  wire result_sign__477;
  wire result_sign__573;
  wire [7:0] result_exp__120;
  wire result_sign__574;
  wire result_sign__675;
  wire [7:0] result_exp__180;
  wire result_sign__676;
  wire result_sign__787;
  wire [7:0] result_exp__240;
  wire result_sign__788;
  wire [22:0] result_fraction__109;
  wire [22:0] result_fraction__111;
  wire [8:0] sum__19;
  wire [22:0] result_fraction__227;
  wire [22:0] result_fraction__226;
  wire [8:0] sum__38;
  wire [22:0] result_fraction__344;
  wire [22:0] result_fraction__343;
  wire [8:0] sum__57;
  wire [22:0] result_fraction__461;
  wire [22:0] result_fraction__460;
  wire [8:0] sum__76;
  wire [22:0] result_fraction__110;
  wire [22:0] nan_fraction__104;
  wire [22:0] result_fraction__112;
  wire [22:0] nan_fraction__103;
  wire [22:0] result_fraction__229;
  wire [22:0] nan_fraction__131;
  wire [22:0] result_fraction__228;
  wire [22:0] nan_fraction__130;
  wire [22:0] result_fraction__346;
  wire [22:0] nan_fraction__160;
  wire [22:0] result_fraction__345;
  wire [22:0] nan_fraction__159;
  wire [22:0] result_fraction__463;
  wire [22:0] nan_fraction__189;
  wire [22:0] result_fraction__462;
  wire [22:0] nan_fraction__188;
  wire [22:0] result_fraction__114;
  wire [22:0] result_fraction__113;
  wire [7:0] y_sq_bexp__1;
  wire [7:0] x_bexp__820;
  wire [22:0] result_fraction__231;
  wire [22:0] result_fraction__230;
  wire [7:0] y_sq_bexp__6;
  wire [7:0] x_bexp__821;
  wire [22:0] result_fraction__348;
  wire [22:0] result_fraction__347;
  wire [7:0] y_sq_bexp__10;
  wire [7:0] x_bexp__822;
  wire [22:0] result_fraction__465;
  wire [22:0] result_fraction__464;
  wire [7:0] y_sq_bexp__14;
  wire [7:0] x_bexp__823;
  wire [22:0] y_sq_fraction;
  wire [7:0] incremented_sum__94;
  wire [22:0] y_sq_fraction__3;
  wire [7:0] incremented_sum__112;
  wire [22:0] y_sq_fraction__6;
  wire [7:0] incremented_sum__130;
  wire [22:0] y_sq_fraction__9;
  wire [7:0] incremented_sum__148;
  wire [27:0] wide_y__37;
  wire [7:0] x_sq_bexpbs_difference__1;
  wire [27:0] wide_y__75;
  wire [7:0] x_sq_bexpbs_difference__2;
  wire [27:0] wide_y__113;
  wire [7:0] x_sq_bexpbs_difference__3;
  wire [27:0] wide_y__151;
  wire [7:0] x_sq_bexpbs_difference__4;
  wire [27:0] wide_y__38;
  wire [7:0] sub_172687;
  wire [27:0] wide_y__76;
  wire [7:0] sub_172689;
  wire [27:0] wide_y__114;
  wire [7:0] sub_172691;
  wire [27:0] wide_y__152;
  wire [7:0] sub_172693;
  wire [27:0] dropped__19;
  wire [27:0] dropped__38;
  wire [27:0] dropped__57;
  wire [27:0] dropped__76;
  wire [7:0] x_sq_bexp__2;
  wire [7:0] x_bexp__824;
  wire [7:0] x_sq_bexp__5;
  wire [7:0] x_bexp__825;
  wire [7:0] x_sq_bexp__10;
  wire [7:0] x_bexp__826;
  wire [7:0] x_sq_bexp__14;
  wire [7:0] x_bexp__827;
  wire [22:0] x_sq_fraction;
  wire [27:0] sticky__59;
  wire [22:0] x_sq_fraction__1;
  wire [27:0] sticky__118;
  wire [22:0] x_sq_fraction__6;
  wire [27:0] sticky__177;
  wire [22:0] x_sq_fraction__9;
  wire [27:0] sticky__236;
  wire [27:0] x_sqddend_y;
  wire [27:0] x_sqddend_y__1;
  wire [27:0] x_sqddend_y__2;
  wire [27:0] x_sqddend_y__3;
  wire [24:0] wide_x__153;
  wire [24:0] wide_x__154;
  wire [24:0] wide_x__155;
  wire [24:0] wide_x__156;
  wire [2:0] bit_slice_172762;
  wire [24:0] carry_fraction__155;
  wire [2:0] bit_slice_172764;
  wire [24:0] carry_fraction__158;
  wire [2:0] bit_slice_172766;
  wire [24:0] carry_fraction__161;
  wire [2:0] bit_slice_172768;
  wire [24:0] carry_fraction__164;
  wire [27:0] concat_172778;
  wire [27:0] concat_172779;
  wire [27:0] concat_172780;
  wire [27:0] concat_172781;
  wire [28:0] one_hot_172782;
  wire [28:0] one_hot_172783;
  wire [28:0] one_hot_172784;
  wire [28:0] one_hot_172785;
  wire [4:0] encode_172786;
  wire [4:0] encode_172787;
  wire [4:0] encode_172788;
  wire [4:0] encode_172789;
  wire cancel__19;
  wire carry_bit__19;
  wire [22:0] result_fraction__536;
  wire cancel__38;
  wire carry_bit__38;
  wire [22:0] result_fraction__603;
  wire cancel__57;
  wire carry_bit__57;
  wire [22:0] result_fraction__670;
  wire cancel__76;
  wire carry_bit__76;
  wire [22:0] result_fraction__749;
  wire [27:0] leading_zeroes__19;
  wire [27:0] leading_zeroes__38;
  wire [27:0] leading_zeroes__57;
  wire [27:0] leading_zeroes__76;
  wire carry_fraction__154;
  wire carry_fraction__153;
  wire [26:0] concat_172839;
  wire [27:0] add_172840;
  wire carry_fraction__157;
  wire carry_fraction__156;
  wire [26:0] concat_172846;
  wire [27:0] add_172847;
  wire carry_fraction__160;
  wire carry_fraction__159;
  wire [26:0] concat_172853;
  wire [27:0] add_172854;
  wire carry_fraction__163;
  wire carry_fraction__162;
  wire [26:0] concat_172860;
  wire [27:0] add_172861;
  wire [2:0] concat_172862;
  wire [26:0] carry_fraction__38;
  wire [26:0] cancel_fraction__19;
  wire [2:0] concat_172865;
  wire [26:0] carry_fraction__76;
  wire [26:0] cancel_fraction__38;
  wire [2:0] concat_172868;
  wire [26:0] carry_fraction__114;
  wire [26:0] cancel_fraction__57;
  wire [2:0] concat_172871;
  wire [26:0] carry_fraction__152;
  wire [26:0] cancel_fraction__76;
  wire [26:0] shifted_fraction__19;
  wire [26:0] shifted_fraction__38;
  wire [26:0] shifted_fraction__57;
  wire [26:0] shifted_fraction__76;
  wire result_sign__1100;
  wire result_sign__1101;
  wire result_sign__1102;
  wire result_sign__1103;
  wire [2:0] normal_chunk__19;
  wire [2:0] fraction_shift__261;
  wire [1:0] half_way_chunk__19;
  wire [2:0] normal_chunk__38;
  wire [2:0] fraction_shift__296;
  wire [1:0] half_way_chunk__38;
  wire [2:0] normal_chunk__57;
  wire [2:0] fraction_shift__331;
  wire [1:0] half_way_chunk__57;
  wire [2:0] normal_chunk__76;
  wire [2:0] fraction_shift__366;
  wire [1:0] half_way_chunk__76;
  wire result_sign__478;
  wire [24:0] add_172913;
  wire result_sign__575;
  wire [24:0] add_172917;
  wire result_sign__677;
  wire [24:0] add_172921;
  wire result_sign__789;
  wire [24:0] add_172925;
  wire do_round_up__39;
  wire do_round_up__78;
  wire do_round_up__117;
  wire do_round_up__156;
  wire [27:0] rounded_fraction__19;
  wire [27:0] rounded_fraction__38;
  wire [27:0] rounded_fraction__57;
  wire [27:0] rounded_fraction__76;
  wire result_sign__479;
  wire [7:0] x_bexp__592;
  wire rounding_carry__19;
  wire result_sign__576;
  wire [7:0] x_bexp__610;
  wire rounding_carry__38;
  wire result_sign__678;
  wire [7:0] x_bexp__628;
  wire rounding_carry__57;
  wire result_sign__790;
  wire [7:0] x_bexp__646;
  wire rounding_carry__76;
  wire result_sign__480;
  wire [8:0] add_172963;
  wire result_sign__577;
  wire [8:0] add_172967;
  wire result_sign__679;
  wire [8:0] add_172971;
  wire result_sign__791;
  wire [8:0] add_172975;
  wire [9:0] add_172998;
  wire [9:0] add_173001;
  wire [9:0] add_173004;
  wire [9:0] add_173007;
  wire [9:0] wide_exponent__55;
  wire [9:0] wide_exponent__112;
  wire [9:0] wide_exponent__169;
  wire [9:0] wide_exponent__226;
  wire [9:0] wide_exponent__56;
  wire [9:0] wide_exponent__113;
  wire [9:0] wide_exponent__170;
  wire [9:0] wide_exponent__227;
  wire [7:0] high_exp__138;
  wire [22:0] result_fraction__537;
  wire [7:0] high_exp__139;
  wire [22:0] result_fraction__538;
  wire [8:0] wide_exponent__57;
  wire [7:0] high_exp__204;
  wire [22:0] result_fraction__604;
  wire [7:0] high_exp__205;
  wire [22:0] result_fraction__605;
  wire [8:0] wide_exponent__114;
  wire [7:0] high_exp__272;
  wire [22:0] result_fraction__671;
  wire [7:0] high_exp__273;
  wire [22:0] result_fraction__672;
  wire [8:0] wide_exponent__171;
  wire [7:0] high_exp__346;
  wire [22:0] result_fraction__750;
  wire [7:0] high_exp__347;
  wire [22:0] result_fraction__751;
  wire [8:0] wide_exponent__228;
  wire eq_173058;
  wire eq_173060;
  wire eq_173063;
  wire eq_173065;
  wire eq_173068;
  wire eq_173070;
  wire eq_173073;
  wire eq_173075;
  wire [22:0] result_fraction__539;
  wire [22:0] result_fraction__540;
  wire [22:0] result_fraction__606;
  wire [22:0] result_fraction__607;
  wire [22:0] result_fraction__673;
  wire [22:0] result_fraction__674;
  wire [22:0] result_fraction__752;
  wire [22:0] result_fraction__753;
  wire [2:0] fraction_shift__384;
  wire [2:0] fraction_shift__262;
  wire is_operand_inf__19;
  wire and_reduce_173112;
  wire [2:0] fraction_shift__402;
  wire [2:0] fraction_shift__297;
  wire is_operand_inf__38;
  wire and_reduce_173120;
  wire [2:0] fraction_shift__420;
  wire [2:0] fraction_shift__332;
  wire is_operand_inf__57;
  wire and_reduce_173128;
  wire [2:0] fraction_shift__438;
  wire [2:0] fraction_shift__367;
  wire is_operand_inf__76;
  wire and_reduce_173136;
  wire [2:0] fraction_shift__57;
  wire [2:0] fraction_shift__114;
  wire [2:0] fraction_shift__171;
  wire [2:0] fraction_shift__228;
  wire is_result_nan__39;
  wire [27:0] shrl_173155;
  wire is_result_nan__78;
  wire [27:0] shrl_173158;
  wire is_result_nan__117;
  wire [27:0] shrl_173161;
  wire is_result_nan__156;
  wire [27:0] shrl_173164;
  wire [7:0] high_exp__140;
  wire [22:0] result_fraction__115;
  wire [7:0] high_exp__206;
  wire [22:0] result_fraction__232;
  wire [7:0] high_exp__274;
  wire [22:0] result_fraction__349;
  wire [7:0] high_exp__348;
  wire [22:0] result_fraction__466;
  wire [7:0] result_exponent__19;
  wire [22:0] result_fraction__116;
  wire [22:0] nan_fraction__105;
  wire [7:0] result_exponent__38;
  wire [22:0] result_fraction__233;
  wire [22:0] nan_fraction__132;
  wire [7:0] result_exponent__57;
  wire [22:0] result_fraction__350;
  wire [22:0] nan_fraction__161;
  wire [7:0] result_exponent__76;
  wire [22:0] result_fraction__467;
  wire [22:0] nan_fraction__190;
  wire [7:0] uexp;
  wire [22:0] result_fraction__117;
  wire result_sign__828;
  wire [7:0] uexp__1;
  wire [22:0] result_fraction__234;
  wire result_sign__829;
  wire [7:0] uexp__2;
  wire [22:0] result_fraction__351;
  wire result_sign__830;
  wire [7:0] uexp__3;
  wire [22:0] result_fraction__468;
  wire result_sign__831;
  wire [24:0] sel_173230;
  wire [24:0] sel_173231;
  wire [24:0] sel_173232;
  wire [24:0] sel_173233;
  wire [6:0] add_173250;
  wire [6:0] add_173251;
  wire [6:0] add_173252;
  wire [6:0] add_173253;
  wire [7:0] add_173276;
  wire [7:0] add_173280;
  wire [7:0] add_173284;
  wire [7:0] add_173288;
  wire ugt_173291;
  wire ugt_173296;
  wire ugt_173301;
  wire ugt_173306;
  wire [31:0] shifting_bit_mask__1;
  wire [28:0] sel_173312;
  wire [31:0] shifting_bit_mask__100;
  wire [28:0] sel_173315;
  wire [31:0] shifting_bit_mask__101;
  wire [28:0] sel_173318;
  wire [31:0] shifting_bit_mask__102;
  wire [28:0] sel_173321;
  wire [31:0] temp__2;
  wire result_sign__832;
  wire [31:0] temp__27;
  wire result_sign__833;
  wire [31:0] temp__52;
  wire result_sign__834;
  wire [31:0] temp__77;
  wire result_sign__835;
  wire [1:0] concat_173339;
  wire [1:0] concat_173344;
  wire [1:0] concat_173349;
  wire [1:0] concat_173354;
  wire ule_173358;
  wire [30:0] sub_173360;
  wire ule_173361;
  wire [30:0] sub_173363;
  wire ule_173364;
  wire [30:0] sub_173366;
  wire ule_173367;
  wire [30:0] sub_173369;
  wire [1:0] sel_173371;
  wire [22:0] result_fraction__888;
  wire [1:0] sel_173375;
  wire [22:0] result_fraction__889;
  wire [1:0] sel_173379;
  wire [22:0] result_fraction__890;
  wire [1:0] sel_173383;
  wire [22:0] result_fraction__891;
  wire [31:0] shifting_bit_mask__2;
  wire [27:0] sel_173388;
  wire [31:0] shifting_bit_mask__103;
  wire [27:0] sel_173391;
  wire [31:0] shifting_bit_mask__104;
  wire [27:0] sel_173394;
  wire [31:0] shifting_bit_mask__105;
  wire [27:0] sel_173397;
  wire [31:0] temp__3;
  wire result_sign__836;
  wire [31:0] temp__28;
  wire result_sign__837;
  wire [31:0] temp__53;
  wire result_sign__838;
  wire [31:0] temp__78;
  wire result_sign__839;
  wire [2:0] concat_173415;
  wire [2:0] concat_173420;
  wire [2:0] concat_173425;
  wire [2:0] concat_173430;
  wire ule_173434;
  wire [30:0] sub_173436;
  wire ule_173437;
  wire [30:0] sub_173439;
  wire ule_173440;
  wire [30:0] sub_173442;
  wire ule_173443;
  wire [30:0] sub_173445;
  wire [2:0] sel_173447;
  wire [2:0] sel_173451;
  wire [2:0] sel_173455;
  wire [2:0] sel_173459;
  wire [31:0] shifting_bit_mask__3;
  wire [26:0] sel_173464;
  wire [31:0] shifting_bit_mask__106;
  wire [26:0] sel_173467;
  wire [31:0] shifting_bit_mask__107;
  wire [26:0] sel_173470;
  wire [31:0] shifting_bit_mask__108;
  wire [26:0] sel_173473;
  wire [31:0] temp__4;
  wire result_sign__840;
  wire [31:0] temp__29;
  wire result_sign__841;
  wire [31:0] temp__54;
  wire result_sign__842;
  wire [31:0] temp__79;
  wire result_sign__843;
  wire [3:0] concat_173491;
  wire [3:0] concat_173496;
  wire [3:0] concat_173501;
  wire [3:0] concat_173506;
  wire ule_173510;
  wire [30:0] sub_173512;
  wire ule_173513;
  wire [30:0] sub_173515;
  wire ule_173516;
  wire [30:0] sub_173518;
  wire ule_173519;
  wire [30:0] sub_173521;
  wire [3:0] sel_173523;
  wire [3:0] sel_173527;
  wire [3:0] sel_173531;
  wire [3:0] sel_173535;
  wire [31:0] shifting_bit_mask__4;
  wire [25:0] sel_173540;
  wire [31:0] shifting_bit_mask__109;
  wire [25:0] sel_173543;
  wire [31:0] shifting_bit_mask__110;
  wire [25:0] sel_173546;
  wire [31:0] shifting_bit_mask__111;
  wire [25:0] sel_173549;
  wire [31:0] temp__5;
  wire result_sign__844;
  wire [31:0] temp__30;
  wire result_sign__845;
  wire [31:0] temp__55;
  wire result_sign__846;
  wire [31:0] temp__80;
  wire result_sign__847;
  wire [4:0] concat_173567;
  wire [4:0] concat_173572;
  wire [4:0] concat_173577;
  wire [4:0] concat_173582;
  wire ule_173586;
  wire [30:0] sub_173588;
  wire ule_173589;
  wire [30:0] sub_173591;
  wire ule_173592;
  wire [30:0] sub_173594;
  wire ule_173595;
  wire [30:0] sub_173597;
  wire [4:0] sel_173599;
  wire [4:0] sel_173603;
  wire [4:0] sel_173607;
  wire [4:0] sel_173611;
  wire [31:0] shifting_bit_mask__5;
  wire [24:0] sel_173616;
  wire [31:0] shifting_bit_mask__112;
  wire [24:0] sel_173619;
  wire [31:0] shifting_bit_mask__113;
  wire [24:0] sel_173622;
  wire [31:0] shifting_bit_mask__114;
  wire [24:0] sel_173625;
  wire [31:0] temp__6;
  wire result_sign__848;
  wire [31:0] temp__31;
  wire result_sign__849;
  wire [31:0] temp__56;
  wire result_sign__850;
  wire [31:0] temp__81;
  wire result_sign__851;
  wire [5:0] concat_173643;
  wire [5:0] concat_173648;
  wire [5:0] concat_173653;
  wire [5:0] concat_173658;
  wire ule_173662;
  wire [30:0] sub_173664;
  wire ule_173665;
  wire [30:0] sub_173667;
  wire ule_173668;
  wire [30:0] sub_173670;
  wire ule_173671;
  wire [30:0] sub_173673;
  wire [5:0] sel_173675;
  wire [5:0] sel_173679;
  wire [5:0] sel_173683;
  wire [5:0] sel_173687;
  wire [31:0] shifting_bit_mask__6;
  wire [23:0] sel_173692;
  wire [31:0] shifting_bit_mask__115;
  wire [23:0] sel_173695;
  wire [31:0] shifting_bit_mask__116;
  wire [23:0] sel_173698;
  wire [31:0] shifting_bit_mask__117;
  wire [23:0] sel_173701;
  wire [31:0] temp__7;
  wire result_sign__852;
  wire [7:0] x_bexp__656;
  wire [31:0] temp__32;
  wire result_sign__853;
  wire [7:0] x_bexp__658;
  wire [31:0] temp__57;
  wire result_sign__854;
  wire [7:0] x_bexp__660;
  wire [31:0] temp__82;
  wire result_sign__855;
  wire [7:0] x_bexp__662;
  wire [6:0] concat_173719;
  wire [6:0] concat_173724;
  wire [6:0] concat_173729;
  wire [6:0] concat_173734;
  wire ule_173738;
  wire [30:0] sub_173740;
  wire ule_173741;
  wire [30:0] sub_173743;
  wire ule_173744;
  wire [30:0] sub_173746;
  wire ule_173747;
  wire [30:0] sub_173749;
  wire [6:0] sel_173751;
  wire [6:0] sel_173755;
  wire [6:0] sel_173759;
  wire [6:0] sel_173763;
  wire [31:0] shifting_bit_mask__7;
  wire [22:0] sel_173768;
  wire [31:0] shifting_bit_mask__118;
  wire [22:0] sel_173771;
  wire [31:0] shifting_bit_mask__119;
  wire [22:0] sel_173774;
  wire [31:0] shifting_bit_mask__120;
  wire [22:0] sel_173777;
  wire [31:0] temp__8;
  wire result_sign__856;
  wire [31:0] temp__33;
  wire result_sign__857;
  wire [31:0] temp__58;
  wire result_sign__858;
  wire [31:0] temp__83;
  wire result_sign__859;
  wire [7:0] concat_173795;
  wire [7:0] concat_173800;
  wire [7:0] concat_173805;
  wire [7:0] concat_173810;
  wire ule_173814;
  wire [30:0] sub_173816;
  wire ule_173817;
  wire [30:0] sub_173819;
  wire ule_173820;
  wire [30:0] sub_173822;
  wire ule_173823;
  wire [30:0] sub_173825;
  wire [7:0] sel_173827;
  wire [7:0] sel_173831;
  wire [7:0] sel_173835;
  wire [7:0] sel_173839;
  wire [31:0] shifting_bit_mask__8;
  wire [21:0] sel_173844;
  wire [31:0] shifting_bit_mask__121;
  wire [21:0] sel_173847;
  wire [31:0] shifting_bit_mask__122;
  wire [21:0] sel_173850;
  wire [31:0] shifting_bit_mask__123;
  wire [21:0] sel_173853;
  wire [31:0] temp__9;
  wire result_sign__860;
  wire [31:0] temp__34;
  wire result_sign__861;
  wire [31:0] temp__59;
  wire result_sign__862;
  wire [31:0] temp__84;
  wire result_sign__863;
  wire [8:0] concat_173871;
  wire [8:0] concat_173876;
  wire [8:0] concat_173881;
  wire [8:0] concat_173886;
  wire ule_173890;
  wire [30:0] sub_173892;
  wire ule_173893;
  wire [30:0] sub_173895;
  wire ule_173896;
  wire [30:0] sub_173898;
  wire ule_173899;
  wire [30:0] sub_173901;
  wire [8:0] sel_173903;
  wire [8:0] sel_173907;
  wire [8:0] sel_173911;
  wire [8:0] sel_173915;
  wire [31:0] shifting_bit_mask__9;
  wire [20:0] sel_173920;
  wire [31:0] shifting_bit_mask__124;
  wire [20:0] sel_173923;
  wire [31:0] shifting_bit_mask__125;
  wire [20:0] sel_173926;
  wire [31:0] shifting_bit_mask__126;
  wire [20:0] sel_173929;
  wire [31:0] temp__10;
  wire result_sign__864;
  wire [31:0] temp__35;
  wire result_sign__865;
  wire [31:0] temp__60;
  wire result_sign__866;
  wire [31:0] temp__85;
  wire result_sign__867;
  wire [9:0] concat_173947;
  wire [9:0] concat_173952;
  wire [9:0] concat_173957;
  wire [9:0] concat_173962;
  wire ule_173966;
  wire [30:0] sub_173968;
  wire ule_173969;
  wire [30:0] sub_173971;
  wire ule_173972;
  wire [30:0] sub_173974;
  wire ule_173975;
  wire [30:0] sub_173977;
  wire [9:0] sel_173979;
  wire [9:0] sel_173983;
  wire [9:0] sel_173987;
  wire [9:0] sel_173991;
  wire [31:0] shifting_bit_mask__10;
  wire [19:0] sel_173996;
  wire [31:0] shifting_bit_mask__127;
  wire [19:0] sel_173999;
  wire [31:0] shifting_bit_mask__128;
  wire [19:0] sel_174002;
  wire [31:0] shifting_bit_mask__129;
  wire [19:0] sel_174005;
  wire [31:0] temp__11;
  wire result_sign__868;
  wire [31:0] temp__36;
  wire result_sign__869;
  wire [31:0] temp__61;
  wire result_sign__870;
  wire [31:0] temp__86;
  wire result_sign__871;
  wire [10:0] concat_174023;
  wire [10:0] concat_174028;
  wire [10:0] concat_174033;
  wire [10:0] concat_174038;
  wire ule_174042;
  wire [30:0] sub_174044;
  wire ule_174045;
  wire [30:0] sub_174047;
  wire ule_174048;
  wire [30:0] sub_174050;
  wire ule_174051;
  wire [30:0] sub_174053;
  wire [10:0] sel_174055;
  wire [10:0] sel_174059;
  wire [10:0] sel_174063;
  wire [10:0] sel_174067;
  wire [31:0] shifting_bit_mask__11;
  wire [18:0] sel_174072;
  wire [31:0] shifting_bit_mask__130;
  wire [18:0] sel_174075;
  wire [31:0] shifting_bit_mask__131;
  wire [18:0] sel_174078;
  wire [31:0] shifting_bit_mask__132;
  wire [18:0] sel_174081;
  wire [31:0] temp__12;
  wire result_sign__792;
  wire result_sign__872;
  wire [31:0] temp__37;
  wire result_sign__793;
  wire result_sign__873;
  wire [31:0] temp__62;
  wire result_sign__794;
  wire result_sign__874;
  wire [31:0] temp__87;
  wire result_sign__795;
  wire result_sign__875;
  wire [11:0] concat_174104;
  wire [11:0] concat_174110;
  wire [11:0] concat_174116;
  wire [11:0] concat_174122;
  wire ule_174126;
  wire result_sign__876;
  wire [30:0] sub_174129;
  wire ule_174130;
  wire result_sign__877;
  wire [30:0] sub_174133;
  wire ule_174134;
  wire result_sign__878;
  wire [30:0] sub_174137;
  wire ule_174138;
  wire result_sign__879;
  wire [30:0] sub_174141;
  wire [11:0] sel_174143;
  wire [11:0] sel_174148;
  wire [11:0] sel_174153;
  wire [11:0] sel_174158;
  wire [31:0] shifting_bit_mask__12;
  wire [18:0] sel_174164;
  wire [31:0] shifting_bit_mask__133;
  wire [18:0] sel_174167;
  wire [31:0] shifting_bit_mask__134;
  wire [18:0] sel_174170;
  wire [31:0] shifting_bit_mask__135;
  wire [18:0] sel_174173;
  wire [31:0] temp__13;
  wire result_sign__880;
  wire [31:0] temp__38;
  wire result_sign__881;
  wire [31:0] temp__63;
  wire result_sign__882;
  wire [31:0] temp__88;
  wire result_sign__883;
  wire [12:0] concat_174196;
  wire [12:0] concat_174202;
  wire [12:0] concat_174208;
  wire [12:0] concat_174214;
  wire ule_174218;
  wire [30:0] sub_174221;
  wire ule_174222;
  wire [30:0] sub_174225;
  wire ule_174226;
  wire [30:0] sub_174229;
  wire ule_174230;
  wire [30:0] sub_174233;
  wire [12:0] sel_174235;
  wire [12:0] sel_174240;
  wire [12:0] sel_174245;
  wire [12:0] sel_174250;
  wire [31:0] shifting_bit_mask__13;
  wire [19:0] sel_174256;
  wire [31:0] shifting_bit_mask__136;
  wire [19:0] sel_174259;
  wire [31:0] shifting_bit_mask__137;
  wire [19:0] sel_174262;
  wire [31:0] shifting_bit_mask__138;
  wire [19:0] sel_174265;
  wire [31:0] temp__14;
  wire result_sign__884;
  wire [31:0] temp__39;
  wire result_sign__885;
  wire [31:0] temp__64;
  wire result_sign__886;
  wire [31:0] temp__89;
  wire result_sign__887;
  wire [13:0] concat_174288;
  wire [13:0] concat_174294;
  wire [13:0] concat_174300;
  wire [13:0] concat_174306;
  wire ule_174310;
  wire [30:0] sub_174313;
  wire ule_174314;
  wire [30:0] sub_174317;
  wire ule_174318;
  wire [30:0] sub_174321;
  wire ule_174322;
  wire [30:0] sub_174325;
  wire [13:0] sel_174327;
  wire [13:0] sel_174332;
  wire [13:0] sel_174337;
  wire [13:0] sel_174342;
  wire [31:0] shifting_bit_mask__14;
  wire [20:0] sel_174348;
  wire [31:0] shifting_bit_mask__139;
  wire [20:0] sel_174351;
  wire [31:0] shifting_bit_mask__140;
  wire [20:0] sel_174354;
  wire [31:0] shifting_bit_mask__141;
  wire [20:0] sel_174357;
  wire [31:0] temp__15;
  wire result_sign__888;
  wire [31:0] temp__40;
  wire result_sign__889;
  wire [31:0] temp__65;
  wire result_sign__890;
  wire [31:0] temp__90;
  wire result_sign__891;
  wire [14:0] concat_174380;
  wire [14:0] concat_174386;
  wire [14:0] concat_174392;
  wire [14:0] concat_174398;
  wire ule_174402;
  wire [30:0] sub_174405;
  wire ule_174406;
  wire [30:0] sub_174409;
  wire ule_174410;
  wire [30:0] sub_174413;
  wire ule_174414;
  wire [30:0] sub_174417;
  wire [14:0] sel_174419;
  wire [14:0] sel_174424;
  wire [14:0] sel_174429;
  wire [14:0] sel_174434;
  wire [31:0] shifting_bit_mask__15;
  wire [21:0] sel_174440;
  wire [31:0] shifting_bit_mask__142;
  wire [21:0] sel_174443;
  wire [31:0] shifting_bit_mask__143;
  wire [21:0] sel_174446;
  wire [31:0] shifting_bit_mask__144;
  wire [21:0] sel_174449;
  wire [31:0] temp__16;
  wire result_sign__892;
  wire [31:0] temp__41;
  wire result_sign__893;
  wire [31:0] temp__66;
  wire result_sign__894;
  wire [31:0] temp__91;
  wire result_sign__895;
  wire [15:0] concat_174472;
  wire [15:0] concat_174478;
  wire [15:0] concat_174484;
  wire [15:0] concat_174490;
  wire ule_174494;
  wire [30:0] sub_174497;
  wire ule_174498;
  wire [30:0] sub_174501;
  wire ule_174502;
  wire [30:0] sub_174505;
  wire ule_174506;
  wire [30:0] sub_174509;
  wire [15:0] sel_174511;
  wire [15:0] sel_174516;
  wire [15:0] sel_174521;
  wire [15:0] sel_174526;
  wire [31:0] shifting_bit_mask__16;
  wire [22:0] sel_174532;
  wire [31:0] shifting_bit_mask__145;
  wire [22:0] sel_174535;
  wire [31:0] shifting_bit_mask__146;
  wire [22:0] sel_174538;
  wire [31:0] shifting_bit_mask__147;
  wire [22:0] sel_174541;
  wire [31:0] temp__17;
  wire result_sign__896;
  wire [31:0] temp__42;
  wire result_sign__897;
  wire [31:0] temp__67;
  wire result_sign__898;
  wire [31:0] temp__92;
  wire result_sign__899;
  wire [16:0] concat_174564;
  wire [16:0] concat_174570;
  wire [16:0] concat_174576;
  wire [16:0] concat_174582;
  wire ule_174586;
  wire [30:0] sub_174589;
  wire ule_174590;
  wire [30:0] sub_174593;
  wire ule_174594;
  wire [30:0] sub_174597;
  wire ule_174598;
  wire [30:0] sub_174601;
  wire [16:0] sel_174603;
  wire [7:0] x_bexp__652;
  wire [16:0] sel_174608;
  wire [7:0] x_bexp__653;
  wire [16:0] sel_174613;
  wire [7:0] x_bexp__654;
  wire [16:0] sel_174618;
  wire [7:0] x_bexp__655;
  wire [31:0] shifting_bit_mask__17;
  wire [23:0] sel_174624;
  wire [31:0] shifting_bit_mask__148;
  wire [23:0] sel_174627;
  wire [31:0] shifting_bit_mask__149;
  wire [23:0] sel_174630;
  wire [31:0] shifting_bit_mask__150;
  wire [23:0] sel_174633;
  wire [31:0] temp__18;
  wire result_sign__900;
  wire [7:0] x_bexp__657;
  wire [31:0] temp__43;
  wire result_sign__901;
  wire [7:0] x_bexp__659;
  wire [31:0] temp__68;
  wire result_sign__902;
  wire [7:0] x_bexp__661;
  wire [31:0] temp__93;
  wire result_sign__903;
  wire [7:0] x_bexp__663;
  wire [17:0] concat_174656;
  wire [17:0] concat_174662;
  wire [17:0] concat_174668;
  wire [17:0] concat_174674;
  wire ule_174678;
  wire [30:0] sub_174681;
  wire ule_174682;
  wire [30:0] sub_174685;
  wire ule_174686;
  wire [30:0] sub_174689;
  wire ule_174690;
  wire [30:0] sub_174693;
  wire [17:0] sel_174695;
  wire [17:0] sel_174700;
  wire [17:0] sel_174705;
  wire [17:0] sel_174710;
  wire [31:0] shifting_bit_mask__18;
  wire [24:0] sel_174716;
  wire [31:0] shifting_bit_mask__151;
  wire [24:0] sel_174719;
  wire [31:0] shifting_bit_mask__152;
  wire [24:0] sel_174722;
  wire [31:0] shifting_bit_mask__153;
  wire [24:0] sel_174725;
  wire [31:0] temp__19;
  wire result_sign__904;
  wire [31:0] temp__44;
  wire result_sign__905;
  wire [31:0] temp__69;
  wire result_sign__906;
  wire [31:0] temp__94;
  wire result_sign__907;
  wire [18:0] concat_174748;
  wire [18:0] concat_174754;
  wire [18:0] concat_174760;
  wire [18:0] concat_174766;
  wire ule_174770;
  wire [30:0] sub_174773;
  wire ule_174774;
  wire [30:0] sub_174777;
  wire ule_174778;
  wire [30:0] sub_174781;
  wire ule_174782;
  wire [30:0] sub_174785;
  wire [18:0] sel_174787;
  wire [18:0] sel_174792;
  wire [18:0] sel_174797;
  wire [18:0] sel_174802;
  wire [31:0] shifting_bit_mask__19;
  wire [25:0] sel_174808;
  wire [31:0] shifting_bit_mask__154;
  wire [25:0] sel_174811;
  wire [31:0] shifting_bit_mask__155;
  wire [25:0] sel_174814;
  wire [31:0] shifting_bit_mask__156;
  wire [25:0] sel_174817;
  wire [31:0] temp__20;
  wire result_sign__908;
  wire [31:0] temp__45;
  wire result_sign__909;
  wire [31:0] temp__70;
  wire result_sign__910;
  wire [31:0] temp__95;
  wire result_sign__911;
  wire [19:0] concat_174840;
  wire [19:0] concat_174846;
  wire [19:0] concat_174852;
  wire [19:0] concat_174858;
  wire ule_174862;
  wire [30:0] sub_174865;
  wire ule_174866;
  wire [30:0] sub_174869;
  wire ule_174870;
  wire [30:0] sub_174873;
  wire ule_174874;
  wire [30:0] sub_174877;
  wire [19:0] sel_174879;
  wire [19:0] sel_174884;
  wire [19:0] sel_174889;
  wire [19:0] sel_174894;
  wire [31:0] shifting_bit_mask__20;
  wire [26:0] sel_174900;
  wire [31:0] shifting_bit_mask__157;
  wire [26:0] sel_174903;
  wire [31:0] shifting_bit_mask__158;
  wire [26:0] sel_174906;
  wire [31:0] shifting_bit_mask__159;
  wire [26:0] sel_174909;
  wire [31:0] temp__21;
  wire result_sign__912;
  wire [31:0] temp__46;
  wire result_sign__913;
  wire [31:0] temp__71;
  wire result_sign__914;
  wire [31:0] temp__96;
  wire result_sign__915;
  wire [20:0] concat_174932;
  wire [20:0] concat_174938;
  wire [20:0] concat_174944;
  wire [20:0] concat_174950;
  wire ule_174954;
  wire [30:0] sub_174957;
  wire ule_174958;
  wire [30:0] sub_174961;
  wire ule_174962;
  wire [30:0] sub_174965;
  wire ule_174966;
  wire [30:0] sub_174969;
  wire [20:0] sel_174971;
  wire [20:0] sel_174976;
  wire [20:0] sel_174981;
  wire [20:0] sel_174986;
  wire [31:0] shifting_bit_mask__21;
  wire [27:0] sel_174992;
  wire [31:0] shifting_bit_mask__160;
  wire [27:0] sel_174995;
  wire [31:0] shifting_bit_mask__161;
  wire [27:0] sel_174998;
  wire [31:0] shifting_bit_mask__162;
  wire [27:0] sel_175001;
  wire [31:0] temp__22;
  wire result_sign__916;
  wire [31:0] temp__47;
  wire result_sign__917;
  wire [31:0] temp__72;
  wire result_sign__918;
  wire [31:0] temp__97;
  wire result_sign__919;
  wire [21:0] concat_175024;
  wire [21:0] concat_175030;
  wire [21:0] concat_175036;
  wire [21:0] concat_175042;
  wire ule_175046;
  wire [30:0] sub_175049;
  wire ule_175050;
  wire [30:0] sub_175053;
  wire ule_175054;
  wire [30:0] sub_175057;
  wire ule_175058;
  wire [30:0] sub_175061;
  wire [21:0] sel_175063;
  wire [21:0] sel_175068;
  wire [21:0] sel_175073;
  wire [21:0] sel_175078;
  wire [31:0] shifting_bit_mask__22;
  wire [28:0] sel_175084;
  wire [31:0] shifting_bit_mask__163;
  wire [28:0] sel_175087;
  wire [31:0] shifting_bit_mask__164;
  wire [28:0] sel_175090;
  wire [31:0] shifting_bit_mask__165;
  wire [28:0] sel_175093;
  wire [31:0] temp__23;
  wire result_sign__920;
  wire [31:0] temp__48;
  wire result_sign__921;
  wire [31:0] temp__73;
  wire result_sign__922;
  wire [31:0] temp__98;
  wire result_sign__923;
  wire [30:0] scaled_fixed_point_x__50;
  wire [22:0] concat_175116;
  wire [30:0] scaled_fixed_point_x__101;
  wire [22:0] concat_175122;
  wire [30:0] scaled_fixed_point_x__155;
  wire [22:0] concat_175128;
  wire [30:0] scaled_fixed_point_x__209;
  wire [22:0] concat_175134;
  wire ule_175138;
  wire [30:0] sub_175141;
  wire ule_175142;
  wire [30:0] sub_175145;
  wire ule_175146;
  wire [30:0] sub_175149;
  wire ule_175150;
  wire [30:0] sub_175153;
  wire [22:0] sel_175155;
  wire [22:0] sel_175160;
  wire [22:0] sel_175165;
  wire [22:0] sel_175170;
  wire [31:0] shifting_bit_mask__23;
  wire [29:0] sel_175176;
  wire result_sign__924;
  wire [31:0] shifting_bit_mask__166;
  wire [29:0] sel_175181;
  wire result_sign__925;
  wire [31:0] shifting_bit_mask__167;
  wire [29:0] sel_175186;
  wire result_sign__926;
  wire [31:0] shifting_bit_mask__168;
  wire [29:0] sel_175191;
  wire result_sign__927;
  wire [31:0] temp__24;
  wire [31:0] scaled_fixed_point_x__53;
  wire [23:0] concat_175196;
  wire [31:0] temp__49;
  wire [31:0] scaled_fixed_point_x__104;
  wire [23:0] concat_175200;
  wire [31:0] temp__74;
  wire [31:0] scaled_fixed_point_x__158;
  wire [23:0] concat_175204;
  wire [31:0] temp__99;
  wire [31:0] scaled_fixed_point_x__212;
  wire [23:0] concat_175208;
  wire ule_175212;
  wire ule_175216;
  wire ule_175220;
  wire ule_175224;
  wire [30:0] concat_175226;
  wire [23:0] sel_175229;
  wire [30:0] concat_175231;
  wire [23:0] sel_175234;
  wire [30:0] concat_175236;
  wire [23:0] sel_175239;
  wire [30:0] concat_175241;
  wire [23:0] sel_175244;
  wire [30:0] sub_175246;
  wire [30:0] sub_175249;
  wire [30:0] sub_175252;
  wire [30:0] sub_175255;
  wire [30:0] scaled_fixed_point_x__54;
  wire [25:0] add_175262;
  wire [30:0] scaled_fixed_point_x__105;
  wire [25:0] add_175267;
  wire [30:0] scaled_fixed_point_x__159;
  wire [25:0] add_175272;
  wire [30:0] scaled_fixed_point_x__213;
  wire [25:0] add_175277;
  wire [5:0] bit_slice_175281;
  wire [5:0] bit_slice_175285;
  wire [5:0] bit_slice_175289;
  wire [5:0] bit_slice_175293;
  wire [24:0] sel_175294;
  wire [24:0] sel_175297;
  wire [24:0] sel_175300;
  wire [24:0] sel_175303;
  wire result_sign__1120;
  wire [6:0] add_175309;
  wire result_sign__1121;
  wire [6:0] add_175314;
  wire result_sign__1122;
  wire [6:0] add_175319;
  wire result_sign__1123;
  wire [6:0] add_175324;
  wire [7:0] high_exp__141;
  wire [22:0] result_fraction__541;
  wire [7:0] high_exp__207;
  wire [22:0] result_fraction__608;
  wire [7:0] high_exp__275;
  wire [22:0] result_fraction__675;
  wire [7:0] high_exp__349;
  wire [22:0] result_fraction__754;
  wire eq_175342;
  wire eq_175343;
  wire [8:0] add_175344;
  wire eq_175345;
  wire eq_175346;
  wire [8:0] add_175347;
  wire eq_175348;
  wire eq_175349;
  wire [8:0] add_175350;
  wire eq_175351;
  wire eq_175352;
  wire [8:0] add_175353;
  wire [22:0] result_fraction__542;
  wire [22:0] result_fraction__609;
  wire [22:0] result_fraction__676;
  wire [22:0] result_fraction__755;
  wire and_175368;
  wire [7:0] x_bexp__828;
  wire and_175374;
  wire [7:0] x_bexp__829;
  wire and_175380;
  wire [7:0] x_bexp__830;
  wire and_175386;
  wire [7:0] x_bexp__831;
  wire and_175390;
  wire [7:0] x_bexp__593;
  wire [7:0] high_exp__142;
  wire [22:0] nan_fraction__106;
  wire ne_175397;
  wire and_175398;
  wire [7:0] x_bexp__611;
  wire [7:0] high_exp__208;
  wire [22:0] nan_fraction__133;
  wire ne_175405;
  wire and_175406;
  wire [7:0] x_bexp__629;
  wire [7:0] high_exp__276;
  wire [22:0] nan_fraction__162;
  wire ne_175413;
  wire and_175414;
  wire [7:0] x_bexp__647;
  wire [7:0] high_exp__350;
  wire [22:0] nan_fraction__191;
  wire ne_175421;
  wire [31:0] pixel_val;
  wire [31:0] pixel_val__1;
  wire [31:0] pixel_val__2;
  wire [31:0] pixel_val__3;
  wire [31:0] array_175531[4];
  assign array_index_157912 = in_img_unflattened[4'h0];
  assign array_index_157913 = in_img_unflattened[4'h1];
  assign array_index_157914 = in_img_unflattened[4'h4];
  assign array_index_157915 = in_img_unflattened[4'h5];
  assign result_sign__389 = 1'h0;
  assign x_bexp__73 = array_index_157912[30:23];
  assign result_sign__482 = 1'h0;
  assign x_bexp__145 = array_index_157913[30:23];
  assign result_sign__579 = 1'h0;
  assign x_bexp__289 = array_index_157914[30:23];
  assign result_sign__681 = 1'h0;
  assign x_bexp__433 = array_index_157915[30:23];
  assign result_sign__390 = 1'h0;
  assign add_157933 = {result_sign__389, x_bexp__73} + 9'h07f;
  assign x_bexp__664 = 8'h00;
  assign result_sign__94 = 1'h0;
  assign x_fraction__73 = array_index_157912[22:0];
  assign result_sign__483 = 1'h0;
  assign add_157938 = {result_sign__482, x_bexp__145} + 9'h07f;
  assign x_bexp__665 = 8'h00;
  assign result_sign__481 = 1'h0;
  assign x_fraction__145 = array_index_157913[22:0];
  assign result_sign__580 = 1'h0;
  assign add_157943 = {result_sign__579, x_bexp__289} + 9'h07f;
  assign x_bexp__666 = 8'h00;
  assign result_sign__578 = 1'h0;
  assign x_fraction__289 = array_index_157914[22:0];
  assign result_sign__682 = 1'h0;
  assign add_157948 = {result_sign__681, x_bexp__433} + 9'h07f;
  assign x_bexp__667 = 8'h00;
  assign result_sign__680 = 1'h0;
  assign x_fraction__433 = array_index_157915[22:0];
  assign ne_157954 = x_bexp__73 != x_bexp__664;
  assign ne_157959 = x_bexp__145 != x_bexp__665;
  assign ne_157964 = x_bexp__289 != x_bexp__666;
  assign ne_157969 = x_bexp__433 != x_bexp__667;
  assign exp__36 = {result_sign__390, add_157933} + 10'h381;
  assign x_fraction__74 = {result_sign__94, x_fraction__73} | 24'h80_0000;
  assign exp__83 = {result_sign__483, add_157938} + 10'h381;
  assign sign_ext_157977 = {10{ne_157959}};
  assign x_fraction__147 = {result_sign__481, x_fraction__145} | 24'h80_0000;
  assign exp__165 = {result_sign__580, add_157943} + 10'h381;
  assign sign_ext_157981 = {10{ne_157964}};
  assign x_fraction__291 = {result_sign__578, x_fraction__289} | 24'h80_0000;
  assign exp__246 = {result_sign__682, add_157948} + 10'h381;
  assign sign_ext_157985 = {10{ne_157969}};
  assign x_fraction__435 = {result_sign__680, x_fraction__433} | 24'h80_0000;
  assign exp__37 = exp__36 & {10{ne_157954}};
  assign x_fraction__75 = x_fraction__74 & {24{ne_157954}};
  assign result_sign__796 = 1'h0;
  assign result_sign__797 = 1'h0;
  assign exp__85 = exp__83 & sign_ext_157977;
  assign x_fraction__149 = x_fraction__147 & {24{ne_157959}};
  assign result_sign__798 = 1'h0;
  assign result_sign__799 = 1'h0;
  assign exp__167 = exp__165 & sign_ext_157981;
  assign x_fraction__293 = x_fraction__291 & {24{ne_157964}};
  assign result_sign__800 = 1'h0;
  assign result_sign__801 = 1'h0;
  assign exp__248 = exp__246 & sign_ext_157985;
  assign x_fraction__437 = x_fraction__435 & {24{ne_157969}};
  assign result_sign__802 = 1'h0;
  assign result_sign__803 = 1'h0;
  assign concat_158012 = {x_fraction__149, result_sign__798};
  assign concat_158013 = {result_sign__799, x_fraction__149};
  assign concat_158015 = {x_fraction__293, result_sign__800};
  assign concat_158016 = {result_sign__801, x_fraction__293};
  assign concat_158018 = {x_fraction__437, result_sign__802};
  assign concat_158019 = {result_sign__803, x_fraction__437};
  assign sel_158020 = $signed(exp__37) <= $signed(10'h000) ? {result_sign__797, x_fraction__75} : {x_fraction__75, result_sign__796};
  assign sel_158021 = $signed(exp__85) <= $signed(10'h000) ? concat_158013 : concat_158012;
  assign sel_158022 = $signed(exp__167) <= $signed(10'h000) ? concat_158016 : concat_158015;
  assign sel_158023 = $signed(exp__248) <= $signed(10'h000) ? concat_158019 : concat_158018;
  assign result_sign__928 = 1'h0;
  assign fraction__86 = sel_158020[23:1];
  assign result_sign__934 = 1'h0;
  assign fraction__190 = sel_158021[23:1];
  assign result_sign__940 = 1'h0;
  assign fraction__369 = sel_158022[23:1];
  assign result_sign__948 = 1'h0;
  assign fraction__548 = sel_158023[23:1];
  assign fraction__87 = {result_sign__928, fraction__86};
  assign fraction__192 = {result_sign__934, fraction__190};
  assign fraction__371 = {result_sign__940, fraction__369};
  assign fraction__550 = {result_sign__948, fraction__548};
  assign do_round_up__18 = sel_158020[0] & sel_158020[1];
  assign add_158049 = fraction__87 + 24'h00_0001;
  assign do_round_up__40 = sel_158021[0] & sel_158021[1];
  assign add_158051 = fraction__192 + 24'h00_0001;
  assign do_round_up__79 = sel_158022[0] & sel_158022[1];
  assign add_158053 = fraction__371 + 24'h00_0001;
  assign do_round_up__118 = sel_158023[0] & sel_158023[1];
  assign add_158055 = fraction__550 + 24'h00_0001;
  assign fraction__88 = do_round_up__18 ? add_158049 : fraction__87;
  assign fraction__194 = do_round_up__40 ? add_158051 : fraction__192;
  assign fraction__373 = do_round_up__79 ? add_158053 : fraction__371;
  assign fraction__552 = do_round_up__118 ? add_158055 : fraction__550;
  assign add_158065 = exp__37 + 10'h001;
  assign add_158067 = exp__85 + 10'h001;
  assign add_158069 = exp__167 + 10'h001;
  assign add_158071 = exp__248 + 10'h001;
  assign exp__39 = fraction__88[23] ? add_158065 : exp__37;
  assign exp__89 = fraction__194[23] ? add_158067 : exp__85;
  assign exp__171 = fraction__373[23] ? add_158069 : exp__167;
  assign exp__253 = fraction__552[23] ? add_158071 : exp__248;
  assign result_exp__27 = exp__39[8:0];
  assign result_exp__61 = exp__89[8:0];
  assign result_exp__121 = exp__171[8:0];
  assign result_exp__181 = exp__253[8:0];
  assign high_exp__9 = 8'hff;
  assign result_fraction__8 = 23'h00_0000;
  assign result_exp__28 = result_exp__27 & {9{$signed(exp__39) > $signed(10'h000)}};
  assign high_exp__143 = 8'hff;
  assign result_fraction__543 = 23'h00_0000;
  assign result_exp__63 = result_exp__61 & {9{$signed(exp__89) > $signed(10'h000)}};
  assign high_exp__209 = 8'hff;
  assign result_fraction__610 = 23'h00_0000;
  assign result_exp__123 = result_exp__121 & {9{$signed(exp__171) > $signed(10'h000)}};
  assign high_exp__277 = 8'hff;
  assign result_fraction__677 = 23'h00_0000;
  assign result_exp__183 = result_exp__181 & {9{$signed(exp__253) > $signed(10'h000)}};
  assign eq_158104 = x_bexp__73 == high_exp__9;
  assign is_result_nan__3 = x_bexp__145 == high_exp__143;
  assign is_result_nan__24 = x_bexp__289 == high_exp__209;
  assign is_result_nan__84 = x_bexp__433 == high_exp__277;
  assign has_inf_arg__9 = eq_158104 & x_fraction__73 == result_fraction__8;
  assign and_reduce_158122 = &result_exp__28[7:0];
  assign is_subnormal__9 = $signed(exp__39) <= $signed(10'h000);
  assign result_fraction__481 = 23'h00_0000;
  assign has_inf_arg__21 = is_result_nan__3 & x_fraction__145 == result_fraction__543;
  assign and_reduce_158127 = &result_exp__63[7:0];
  assign is_subnormal__21 = $signed(exp__89) <= $signed(10'h000);
  assign result_fraction__544 = 23'h00_0000;
  assign has_inf_arg__41 = is_result_nan__24 & x_fraction__289 == result_fraction__610;
  assign and_reduce_158132 = &result_exp__123[7:0];
  assign is_subnormal__41 = $signed(exp__171) <= $signed(10'h000);
  assign result_fraction__611 = 23'h00_0000;
  assign has_inf_arg__61 = is_result_nan__84 & x_fraction__433 == result_fraction__677;
  assign and_reduce_158137 = &result_exp__183[7:0];
  assign is_subnormal__61 = $signed(exp__253) <= $signed(10'h000);
  assign result_fraction__678 = 23'h00_0000;
  assign ne_158141 = x_fraction__73 != result_fraction__481;
  assign ne_158143 = x_fraction__145 != result_fraction__544;
  assign ne_158145 = x_fraction__289 != result_fraction__611;
  assign ne_158147 = x_fraction__433 != result_fraction__678;
  assign is_result_nan__18 = eq_158104 & ne_158141;
  assign is_result_nan__40 = is_result_nan__3 & ne_158143;
  assign is_result_nan__79 = is_result_nan__24 & ne_158145;
  assign is_result_nan__118 = is_result_nan__84 & ne_158147;
  assign result_fraction__54 = fraction__88[22:0];
  assign or_158158 = is_result_nan__18 | has_inf_arg__9 | result_exp__28[8] | and_reduce_158122;
  assign high_exp__81 = 8'hff;
  assign result_fraction__118 = fraction__194[22:0];
  assign or_158162 = is_result_nan__40 | has_inf_arg__21 | result_exp__63[8] | and_reduce_158127;
  assign high_exp__144 = 8'hff;
  assign result_fraction__235 = fraction__373[22:0];
  assign or_158166 = is_result_nan__79 | has_inf_arg__41 | result_exp__123[8] | and_reduce_158132;
  assign high_exp__210 = 8'hff;
  assign result_fraction__352 = fraction__552[22:0];
  assign or_158170 = is_result_nan__118 | has_inf_arg__61 | result_exp__183[8] | and_reduce_158137;
  assign high_exp__278 = 8'hff;
  assign result_fraction__55 = result_fraction__54 & {23{~(has_inf_arg__9 | result_exp__28[8] | and_reduce_158122 | is_subnormal__9)}};
  assign nan_fraction__9 = 23'h40_0000;
  assign result_exp__29 = or_158158 ? high_exp__81 : result_exp__28[7:0];
  assign x_bexp__668 = 8'h00;
  assign result_fraction__120 = result_fraction__118 & {23{~(has_inf_arg__21 | result_exp__63[8] | and_reduce_158127 | is_subnormal__21)}};
  assign nan_fraction__107 = 23'h40_0000;
  assign result_exp__65 = or_158162 ? high_exp__144 : result_exp__63[7:0];
  assign x_bexp__669 = 8'h00;
  assign result_fraction__237 = result_fraction__235 & {23{~(has_inf_arg__41 | result_exp__123[8] | and_reduce_158132 | is_subnormal__41)}};
  assign nan_fraction__134 = 23'h40_0000;
  assign result_exp__125 = or_158166 ? high_exp__210 : result_exp__123[7:0];
  assign x_bexp__670 = 8'h00;
  assign result_fraction__354 = result_fraction__352 & {23{~(has_inf_arg__61 | result_exp__183[8] | and_reduce_158137 | is_subnormal__61)}};
  assign nan_fraction__163 = 23'h40_0000;
  assign result_exp__185 = or_158170 ? high_exp__278 : result_exp__183[7:0];
  assign x_bexp__671 = 8'h00;
  assign result_fraction__56 = is_result_nan__18 ? nan_fraction__9 : result_fraction__55;
  assign result_fraction__122 = is_result_nan__40 ? nan_fraction__107 : result_fraction__120;
  assign result_fraction__239 = is_result_nan__79 ? nan_fraction__134 : result_fraction__237;
  assign result_fraction__356 = is_result_nan__118 ? nan_fraction__163 : result_fraction__354;
  assign wide_x__18 = {2'h1, result_fraction__56, 3'h0};
  assign wide_x__39 = {2'h1, result_fraction__122, 3'h0};
  assign wide_x__77 = {2'h1, result_fraction__239, 3'h0};
  assign wide_x__115 = {2'h1, result_fraction__356, 3'h0};
  assign x_sign__19 = array_index_157912[31:31];
  assign wide_x__19 = wide_x__18 & {28{result_exp__29 != x_bexp__668}};
  assign x_sign__37 = array_index_157913[31:31];
  assign wide_x__41 = wide_x__39 & {28{result_exp__65 != x_bexp__669}};
  assign x_sign__73 = array_index_157914[31:31];
  assign wide_x__79 = wide_x__77 & {28{result_exp__125 != x_bexp__670}};
  assign x_sign__109 = array_index_157915[31:31];
  assign wide_x__117 = wide_x__115 & {28{result_exp__185 != x_bexp__671}};
  assign result_sign__45 = ~x_sign__19;
  assign neg_158222 = -wide_x__19;
  assign result_sign__98 = ~x_sign__37;
  assign neg_158225 = -wide_x__41;
  assign result_sign__195 = ~x_sign__73;
  assign neg_158228 = -wide_x__79;
  assign result_sign__292 = ~x_sign__109;
  assign neg_158231 = -wide_x__117;
  assign result_sign__46 = ~(eq_158104 & ne_158141) & result_sign__45;
  assign result_sign__100 = ~(is_result_nan__3 & ne_158143) & result_sign__98;
  assign result_sign__197 = ~(is_result_nan__24 & ne_158145) & result_sign__195;
  assign result_sign__294 = ~(is_result_nan__84 & ne_158147) & result_sign__292;
  assign sel_158244 = result_sign__46 ? neg_158222[27:3] : wide_x__19[27:3];
  assign sel_158246 = result_sign__100 ? neg_158225[27:3] : wide_x__41[27:3];
  assign sel_158248 = result_sign__197 ? neg_158228[27:3] : wide_x__79[27:3];
  assign sel_158250 = result_sign__294 ? neg_158231[27:3] : wide_x__117[27:3];
  assign xddend_x__10 = {sel_158244, 3'h0};
  assign xddend_x__19 = {sel_158246, 3'h0};
  assign xddend_x__37 = {sel_158248, 3'h0};
  assign xddend_x__55 = {sel_158250, 3'h0};
  assign fraction__89 = {{1{xddend_x__10[27]}}, xddend_x__10};
  assign neg_158257 = -xddend_x__10;
  assign fraction__196 = {{1{xddend_x__19[27]}}, xddend_x__19};
  assign neg_158259 = -xddend_x__19;
  assign fraction__375 = {{1{xddend_x__37[27]}}, xddend_x__37};
  assign neg_158261 = -xddend_x__37;
  assign fraction__554 = {{1{xddend_x__55[27]}}, xddend_x__55};
  assign neg_158263 = -xddend_x__55;
  assign result_sign__47 = fraction__89[28];
  assign result_sign__102 = fraction__196[28];
  assign result_sign__199 = fraction__375[28];
  assign result_sign__296 = fraction__554[28];
  assign sel_158272 = result_sign__47 ? neg_158257[27:3] : sel_158244;
  assign sel_158273 = result_sign__102 ? neg_158259[27:3] : sel_158246;
  assign sel_158274 = result_sign__199 ? neg_158261[27:3] : sel_158248;
  assign sel_158275 = result_sign__296 ? neg_158263[27:3] : sel_158250;
  assign concat_158284 = {3'h0, {sel_158272[0], sel_158272[1], sel_158272[2], sel_158272[3], sel_158272[4], sel_158272[5], sel_158272[6], sel_158272[7], sel_158272[8], sel_158272[9], sel_158272[10], sel_158272[11], sel_158272[12], sel_158272[13], sel_158272[14], sel_158272[15], sel_158272[16], sel_158272[17], sel_158272[18], sel_158272[19], sel_158272[20], sel_158272[21], sel_158272[22], sel_158272[23], sel_158272[24]}};
  assign concat_158285 = {3'h0, {sel_158273[0], sel_158273[1], sel_158273[2], sel_158273[3], sel_158273[4], sel_158273[5], sel_158273[6], sel_158273[7], sel_158273[8], sel_158273[9], sel_158273[10], sel_158273[11], sel_158273[12], sel_158273[13], sel_158273[14], sel_158273[15], sel_158273[16], sel_158273[17], sel_158273[18], sel_158273[19], sel_158273[20], sel_158273[21], sel_158273[22], sel_158273[23], sel_158273[24]}};
  assign concat_158286 = {3'h0, {sel_158274[0], sel_158274[1], sel_158274[2], sel_158274[3], sel_158274[4], sel_158274[5], sel_158274[6], sel_158274[7], sel_158274[8], sel_158274[9], sel_158274[10], sel_158274[11], sel_158274[12], sel_158274[13], sel_158274[14], sel_158274[15], sel_158274[16], sel_158274[17], sel_158274[18], sel_158274[19], sel_158274[20], sel_158274[21], sel_158274[22], sel_158274[23], sel_158274[24]}};
  assign concat_158287 = {3'h0, {sel_158275[0], sel_158275[1], sel_158275[2], sel_158275[3], sel_158275[4], sel_158275[5], sel_158275[6], sel_158275[7], sel_158275[8], sel_158275[9], sel_158275[10], sel_158275[11], sel_158275[12], sel_158275[13], sel_158275[14], sel_158275[15], sel_158275[16], sel_158275[17], sel_158275[18], sel_158275[19], sel_158275[20], sel_158275[21], sel_158275[22], sel_158275[23], sel_158275[24]}};
  assign one_hot_158288 = {concat_158284[27:0] == 28'h000_0000, concat_158284[27] && concat_158284[26:0] == 27'h000_0000, concat_158284[26] && concat_158284[25:0] == 26'h000_0000, concat_158284[25] && concat_158284[24:0] == 25'h000_0000, concat_158284[24] && concat_158284[23:0] == 24'h00_0000, concat_158284[23] && concat_158284[22:0] == 23'h00_0000, concat_158284[22] && concat_158284[21:0] == 22'h00_0000, concat_158284[21] && concat_158284[20:0] == 21'h00_0000, concat_158284[20] && concat_158284[19:0] == 20'h0_0000, concat_158284[19] && concat_158284[18:0] == 19'h0_0000, concat_158284[18] && concat_158284[17:0] == 18'h0_0000, concat_158284[17] && concat_158284[16:0] == 17'h0_0000, concat_158284[16] && concat_158284[15:0] == 16'h0000, concat_158284[15] && concat_158284[14:0] == 15'h0000, concat_158284[14] && concat_158284[13:0] == 14'h0000, concat_158284[13] && concat_158284[12:0] == 13'h0000, concat_158284[12] && concat_158284[11:0] == 12'h000, concat_158284[11] && concat_158284[10:0] == 11'h000, concat_158284[10] && concat_158284[9:0] == 10'h000, concat_158284[9] && concat_158284[8:0] == 9'h000, concat_158284[8] && concat_158284[7:0] == 8'h00, concat_158284[7] && concat_158284[6:0] == 7'h00, concat_158284[6] && concat_158284[5:0] == 6'h00, concat_158284[5] && concat_158284[4:0] == 5'h00, concat_158284[4] && concat_158284[3:0] == 4'h0, concat_158284[3] && concat_158284[2:0] == 3'h0, concat_158284[2] && concat_158284[1:0] == 2'h0, concat_158284[1] && !concat_158284[0], concat_158284[0]};
  assign one_hot_158289 = {concat_158285[27:0] == 28'h000_0000, concat_158285[27] && concat_158285[26:0] == 27'h000_0000, concat_158285[26] && concat_158285[25:0] == 26'h000_0000, concat_158285[25] && concat_158285[24:0] == 25'h000_0000, concat_158285[24] && concat_158285[23:0] == 24'h00_0000, concat_158285[23] && concat_158285[22:0] == 23'h00_0000, concat_158285[22] && concat_158285[21:0] == 22'h00_0000, concat_158285[21] && concat_158285[20:0] == 21'h00_0000, concat_158285[20] && concat_158285[19:0] == 20'h0_0000, concat_158285[19] && concat_158285[18:0] == 19'h0_0000, concat_158285[18] && concat_158285[17:0] == 18'h0_0000, concat_158285[17] && concat_158285[16:0] == 17'h0_0000, concat_158285[16] && concat_158285[15:0] == 16'h0000, concat_158285[15] && concat_158285[14:0] == 15'h0000, concat_158285[14] && concat_158285[13:0] == 14'h0000, concat_158285[13] && concat_158285[12:0] == 13'h0000, concat_158285[12] && concat_158285[11:0] == 12'h000, concat_158285[11] && concat_158285[10:0] == 11'h000, concat_158285[10] && concat_158285[9:0] == 10'h000, concat_158285[9] && concat_158285[8:0] == 9'h000, concat_158285[8] && concat_158285[7:0] == 8'h00, concat_158285[7] && concat_158285[6:0] == 7'h00, concat_158285[6] && concat_158285[5:0] == 6'h00, concat_158285[5] && concat_158285[4:0] == 5'h00, concat_158285[4] && concat_158285[3:0] == 4'h0, concat_158285[3] && concat_158285[2:0] == 3'h0, concat_158285[2] && concat_158285[1:0] == 2'h0, concat_158285[1] && !concat_158285[0], concat_158285[0]};
  assign one_hot_158290 = {concat_158286[27:0] == 28'h000_0000, concat_158286[27] && concat_158286[26:0] == 27'h000_0000, concat_158286[26] && concat_158286[25:0] == 26'h000_0000, concat_158286[25] && concat_158286[24:0] == 25'h000_0000, concat_158286[24] && concat_158286[23:0] == 24'h00_0000, concat_158286[23] && concat_158286[22:0] == 23'h00_0000, concat_158286[22] && concat_158286[21:0] == 22'h00_0000, concat_158286[21] && concat_158286[20:0] == 21'h00_0000, concat_158286[20] && concat_158286[19:0] == 20'h0_0000, concat_158286[19] && concat_158286[18:0] == 19'h0_0000, concat_158286[18] && concat_158286[17:0] == 18'h0_0000, concat_158286[17] && concat_158286[16:0] == 17'h0_0000, concat_158286[16] && concat_158286[15:0] == 16'h0000, concat_158286[15] && concat_158286[14:0] == 15'h0000, concat_158286[14] && concat_158286[13:0] == 14'h0000, concat_158286[13] && concat_158286[12:0] == 13'h0000, concat_158286[12] && concat_158286[11:0] == 12'h000, concat_158286[11] && concat_158286[10:0] == 11'h000, concat_158286[10] && concat_158286[9:0] == 10'h000, concat_158286[9] && concat_158286[8:0] == 9'h000, concat_158286[8] && concat_158286[7:0] == 8'h00, concat_158286[7] && concat_158286[6:0] == 7'h00, concat_158286[6] && concat_158286[5:0] == 6'h00, concat_158286[5] && concat_158286[4:0] == 5'h00, concat_158286[4] && concat_158286[3:0] == 4'h0, concat_158286[3] && concat_158286[2:0] == 3'h0, concat_158286[2] && concat_158286[1:0] == 2'h0, concat_158286[1] && !concat_158286[0], concat_158286[0]};
  assign one_hot_158291 = {concat_158287[27:0] == 28'h000_0000, concat_158287[27] && concat_158287[26:0] == 27'h000_0000, concat_158287[26] && concat_158287[25:0] == 26'h000_0000, concat_158287[25] && concat_158287[24:0] == 25'h000_0000, concat_158287[24] && concat_158287[23:0] == 24'h00_0000, concat_158287[23] && concat_158287[22:0] == 23'h00_0000, concat_158287[22] && concat_158287[21:0] == 22'h00_0000, concat_158287[21] && concat_158287[20:0] == 21'h00_0000, concat_158287[20] && concat_158287[19:0] == 20'h0_0000, concat_158287[19] && concat_158287[18:0] == 19'h0_0000, concat_158287[18] && concat_158287[17:0] == 18'h0_0000, concat_158287[17] && concat_158287[16:0] == 17'h0_0000, concat_158287[16] && concat_158287[15:0] == 16'h0000, concat_158287[15] && concat_158287[14:0] == 15'h0000, concat_158287[14] && concat_158287[13:0] == 14'h0000, concat_158287[13] && concat_158287[12:0] == 13'h0000, concat_158287[12] && concat_158287[11:0] == 12'h000, concat_158287[11] && concat_158287[10:0] == 11'h000, concat_158287[10] && concat_158287[9:0] == 10'h000, concat_158287[9] && concat_158287[8:0] == 9'h000, concat_158287[8] && concat_158287[7:0] == 8'h00, concat_158287[7] && concat_158287[6:0] == 7'h00, concat_158287[6] && concat_158287[5:0] == 6'h00, concat_158287[5] && concat_158287[4:0] == 5'h00, concat_158287[4] && concat_158287[3:0] == 4'h0, concat_158287[3] && concat_158287[2:0] == 3'h0, concat_158287[2] && concat_158287[1:0] == 2'h0, concat_158287[1] && !concat_158287[0], concat_158287[0]};
  assign encode_158292 = {one_hot_158288[16] | one_hot_158288[17] | one_hot_158288[18] | one_hot_158288[19] | one_hot_158288[20] | one_hot_158288[21] | one_hot_158288[22] | one_hot_158288[23] | one_hot_158288[24] | one_hot_158288[25] | one_hot_158288[26] | one_hot_158288[27] | one_hot_158288[28], one_hot_158288[8] | one_hot_158288[9] | one_hot_158288[10] | one_hot_158288[11] | one_hot_158288[12] | one_hot_158288[13] | one_hot_158288[14] | one_hot_158288[15] | one_hot_158288[24] | one_hot_158288[25] | one_hot_158288[26] | one_hot_158288[27] | one_hot_158288[28], one_hot_158288[4] | one_hot_158288[5] | one_hot_158288[6] | one_hot_158288[7] | one_hot_158288[12] | one_hot_158288[13] | one_hot_158288[14] | one_hot_158288[15] | one_hot_158288[20] | one_hot_158288[21] | one_hot_158288[22] | one_hot_158288[23] | one_hot_158288[28], one_hot_158288[2] | one_hot_158288[3] | one_hot_158288[6] | one_hot_158288[7] | one_hot_158288[10] | one_hot_158288[11] | one_hot_158288[14] | one_hot_158288[15] | one_hot_158288[18] | one_hot_158288[19] | one_hot_158288[22] | one_hot_158288[23] | one_hot_158288[26] | one_hot_158288[27], one_hot_158288[1] | one_hot_158288[3] | one_hot_158288[5] | one_hot_158288[7] | one_hot_158288[9] | one_hot_158288[11] | one_hot_158288[13] | one_hot_158288[15] | one_hot_158288[17] | one_hot_158288[19] | one_hot_158288[21] | one_hot_158288[23] | one_hot_158288[25] | one_hot_158288[27]};
  assign encode_158293 = {one_hot_158289[16] | one_hot_158289[17] | one_hot_158289[18] | one_hot_158289[19] | one_hot_158289[20] | one_hot_158289[21] | one_hot_158289[22] | one_hot_158289[23] | one_hot_158289[24] | one_hot_158289[25] | one_hot_158289[26] | one_hot_158289[27] | one_hot_158289[28], one_hot_158289[8] | one_hot_158289[9] | one_hot_158289[10] | one_hot_158289[11] | one_hot_158289[12] | one_hot_158289[13] | one_hot_158289[14] | one_hot_158289[15] | one_hot_158289[24] | one_hot_158289[25] | one_hot_158289[26] | one_hot_158289[27] | one_hot_158289[28], one_hot_158289[4] | one_hot_158289[5] | one_hot_158289[6] | one_hot_158289[7] | one_hot_158289[12] | one_hot_158289[13] | one_hot_158289[14] | one_hot_158289[15] | one_hot_158289[20] | one_hot_158289[21] | one_hot_158289[22] | one_hot_158289[23] | one_hot_158289[28], one_hot_158289[2] | one_hot_158289[3] | one_hot_158289[6] | one_hot_158289[7] | one_hot_158289[10] | one_hot_158289[11] | one_hot_158289[14] | one_hot_158289[15] | one_hot_158289[18] | one_hot_158289[19] | one_hot_158289[22] | one_hot_158289[23] | one_hot_158289[26] | one_hot_158289[27], one_hot_158289[1] | one_hot_158289[3] | one_hot_158289[5] | one_hot_158289[7] | one_hot_158289[9] | one_hot_158289[11] | one_hot_158289[13] | one_hot_158289[15] | one_hot_158289[17] | one_hot_158289[19] | one_hot_158289[21] | one_hot_158289[23] | one_hot_158289[25] | one_hot_158289[27]};
  assign encode_158294 = {one_hot_158290[16] | one_hot_158290[17] | one_hot_158290[18] | one_hot_158290[19] | one_hot_158290[20] | one_hot_158290[21] | one_hot_158290[22] | one_hot_158290[23] | one_hot_158290[24] | one_hot_158290[25] | one_hot_158290[26] | one_hot_158290[27] | one_hot_158290[28], one_hot_158290[8] | one_hot_158290[9] | one_hot_158290[10] | one_hot_158290[11] | one_hot_158290[12] | one_hot_158290[13] | one_hot_158290[14] | one_hot_158290[15] | one_hot_158290[24] | one_hot_158290[25] | one_hot_158290[26] | one_hot_158290[27] | one_hot_158290[28], one_hot_158290[4] | one_hot_158290[5] | one_hot_158290[6] | one_hot_158290[7] | one_hot_158290[12] | one_hot_158290[13] | one_hot_158290[14] | one_hot_158290[15] | one_hot_158290[20] | one_hot_158290[21] | one_hot_158290[22] | one_hot_158290[23] | one_hot_158290[28], one_hot_158290[2] | one_hot_158290[3] | one_hot_158290[6] | one_hot_158290[7] | one_hot_158290[10] | one_hot_158290[11] | one_hot_158290[14] | one_hot_158290[15] | one_hot_158290[18] | one_hot_158290[19] | one_hot_158290[22] | one_hot_158290[23] | one_hot_158290[26] | one_hot_158290[27], one_hot_158290[1] | one_hot_158290[3] | one_hot_158290[5] | one_hot_158290[7] | one_hot_158290[9] | one_hot_158290[11] | one_hot_158290[13] | one_hot_158290[15] | one_hot_158290[17] | one_hot_158290[19] | one_hot_158290[21] | one_hot_158290[23] | one_hot_158290[25] | one_hot_158290[27]};
  assign encode_158295 = {one_hot_158291[16] | one_hot_158291[17] | one_hot_158291[18] | one_hot_158291[19] | one_hot_158291[20] | one_hot_158291[21] | one_hot_158291[22] | one_hot_158291[23] | one_hot_158291[24] | one_hot_158291[25] | one_hot_158291[26] | one_hot_158291[27] | one_hot_158291[28], one_hot_158291[8] | one_hot_158291[9] | one_hot_158291[10] | one_hot_158291[11] | one_hot_158291[12] | one_hot_158291[13] | one_hot_158291[14] | one_hot_158291[15] | one_hot_158291[24] | one_hot_158291[25] | one_hot_158291[26] | one_hot_158291[27] | one_hot_158291[28], one_hot_158291[4] | one_hot_158291[5] | one_hot_158291[6] | one_hot_158291[7] | one_hot_158291[12] | one_hot_158291[13] | one_hot_158291[14] | one_hot_158291[15] | one_hot_158291[20] | one_hot_158291[21] | one_hot_158291[22] | one_hot_158291[23] | one_hot_158291[28], one_hot_158291[2] | one_hot_158291[3] | one_hot_158291[6] | one_hot_158291[7] | one_hot_158291[10] | one_hot_158291[11] | one_hot_158291[14] | one_hot_158291[15] | one_hot_158291[18] | one_hot_158291[19] | one_hot_158291[22] | one_hot_158291[23] | one_hot_158291[26] | one_hot_158291[27], one_hot_158291[1] | one_hot_158291[3] | one_hot_158291[5] | one_hot_158291[7] | one_hot_158291[9] | one_hot_158291[11] | one_hot_158291[13] | one_hot_158291[15] | one_hot_158291[17] | one_hot_158291[19] | one_hot_158291[21] | one_hot_158291[23] | one_hot_158291[25] | one_hot_158291[27]};
  assign result_fraction__482 = 23'h00_0000;
  assign result_fraction__545 = 23'h00_0000;
  assign result_fraction__612 = 23'h00_0000;
  assign result_fraction__679 = 23'h00_0000;
  assign cancel__10 = |encode_158292[4:1];
  assign carry_bit__9 = sel_158272[24];
  assign leading_zeroes__9 = {result_fraction__482, encode_158292};
  assign cancel__20 = |encode_158293[4:1];
  assign carry_bit__20 = sel_158273[24];
  assign leading_zeroes__20 = {result_fraction__545, encode_158293};
  assign array_index_158318 = in_img_unflattened[4'h2];
  assign cancel__39 = |encode_158294[4:1];
  assign carry_bit__39 = sel_158274[24];
  assign leading_zeroes__39 = {result_fraction__612, encode_158294};
  assign cancel__58 = |encode_158295[4:1];
  assign carry_bit__58 = sel_158275[24];
  assign leading_zeroes__58 = {result_fraction__679, encode_158295};
  assign array_index_158331 = in_img_unflattened[4'h6];
  assign add_158335 = leading_zeroes__9 + 28'hfff_ffff;
  assign add_158339 = leading_zeroes__20 + 28'hfff_ffff;
  assign x_bexp__157 = array_index_158318[30:23];
  assign add_158344 = leading_zeroes__39 + 28'hfff_ffff;
  assign add_158348 = leading_zeroes__58 + 28'hfff_ffff;
  assign x_bexp__445 = array_index_158331[30:23];
  assign cancel_fraction__9 = add_158335 >= 28'h000_001b ? 27'h000_0000 : {sel_158272[23:0], 3'h0} << add_158335;
  assign result_sign__956 = 1'h0;
  assign cancel_fraction__20 = add_158339 >= 28'h000_001b ? 27'h000_0000 : {sel_158273[23:0], 3'h0} << add_158339;
  assign result_sign__957 = 1'h0;
  assign cancel_fraction__39 = add_158344 >= 28'h000_001b ? 27'h000_0000 : {sel_158274[23:0], 3'h0} << add_158344;
  assign result_sign__958 = 1'h0;
  assign cancel_fraction__58 = add_158348 >= 28'h000_001b ? 27'h000_0000 : {sel_158275[23:0], 3'h0} << add_158348;
  assign result_sign__959 = 1'h0;
  assign concat_158374 = {~(carry_bit__9 | cancel__10), ~(carry_bit__9 | ~cancel__10), ~(~carry_bit__9 | cancel__10)};
  assign concat_158379 = {~(carry_bit__20 | cancel__20), ~(carry_bit__20 | ~cancel__20), ~(~carry_bit__20 | cancel__20)};
  assign concat_158384 = {~(carry_bit__39 | cancel__39), ~(carry_bit__39 | ~cancel__39), ~(~carry_bit__39 | cancel__39)};
  assign concat_158389 = {~(carry_bit__58 | cancel__58), ~(carry_bit__58 | ~cancel__58), ~(~carry_bit__58 | cancel__58)};
  assign result_sign__960 = 1'h0;
  assign one_hot_sel_158396 = sel_158272[24:1] & {24{concat_158374[0]}} | cancel_fraction__9[26:3] & {24{concat_158374[1]}} | sel_158272[23:0] & {24{concat_158374[2]}};
  assign result_sign__1104 = 1'h0;
  assign add_158398 = {result_sign__956, x_bexp__145[7]} + 2'h1;
  assign result_sign__961 = 1'h0;
  assign one_hot_sel_158402 = sel_158273[24:1] & {24{concat_158379[0]}} | cancel_fraction__20[26:3] & {24{concat_158379[1]}} | sel_158273[23:0] & {24{concat_158379[2]}};
  assign result_sign__1106 = 1'h0;
  assign add_158404 = {result_sign__957, x_bexp__157[7]} + 2'h1;
  assign x_bexp__672 = 8'h00;
  assign result_sign__484 = 1'h0;
  assign x_fraction__157 = array_index_158318[22:0];
  assign result_sign__962 = 1'h0;
  assign one_hot_sel_158411 = sel_158274[24:1] & {24{concat_158384[0]}} | cancel_fraction__39[26:3] & {24{concat_158384[1]}} | sel_158274[23:0] & {24{concat_158384[2]}};
  assign result_sign__1108 = 1'h0;
  assign add_158413 = {result_sign__958, x_bexp__433[7]} + 2'h1;
  assign result_sign__963 = 1'h0;
  assign one_hot_sel_158417 = sel_158275[24:1] & {24{concat_158389[0]}} | cancel_fraction__58[26:3] & {24{concat_158389[1]}} | sel_158275[23:0] & {24{concat_158389[2]}};
  assign result_sign__1112 = 1'h0;
  assign add_158419 = {result_sign__959, x_bexp__445[7]} + 2'h1;
  assign x_bexp__673 = 8'h00;
  assign result_sign__683 = 1'h0;
  assign x_fraction__445 = array_index_158331[22:0];
  assign ne_158434 = x_bexp__157 != x_bexp__672;
  assign ne_158447 = x_bexp__445 != x_bexp__673;
  assign nor_158451 = ~(~carry_bit__9 | cancel__10 | ~sel_158272[0]);
  assign result_sign__1116 = 1'h0;
  assign add_158453 = {result_sign__960, one_hot_sel_158396} + 25'h000_0001;
  assign exp__40 = {result_sign__1104, add_158398, x_bexp__145[6:0]} + 10'h381;
  assign nor_158456 = ~(~carry_bit__20 | cancel__20 | ~sel_158273[0]);
  assign result_sign__1117 = 1'h0;
  assign add_158458 = {result_sign__961, one_hot_sel_158402} + 25'h000_0001;
  assign exp__91 = {result_sign__1106, add_158404, x_bexp__157[6:0]} + 10'h381;
  assign sign_ext_158460 = {10{ne_158434}};
  assign x_fraction__159 = {result_sign__484, x_fraction__157} | 24'h80_0000;
  assign nor_158464 = ~(~carry_bit__39 | cancel__39 | ~sel_158274[0]);
  assign result_sign__1118 = 1'h0;
  assign add_158466 = {result_sign__962, one_hot_sel_158411} + 25'h000_0001;
  assign exp__173 = {result_sign__1108, add_158413, x_bexp__433[6:0]} + 10'h381;
  assign nor_158469 = ~(~carry_bit__58 | cancel__58 | ~sel_158275[0]);
  assign result_sign__1119 = 1'h0;
  assign add_158471 = {result_sign__963, one_hot_sel_158417} + 25'h000_0001;
  assign exp__255 = {result_sign__1112, add_158419, x_bexp__445[6:0]} + 10'h381;
  assign sign_ext_158473 = {10{ne_158447}};
  assign x_fraction__447 = {result_sign__683, x_fraction__445} | 24'h80_0000;
  assign do_round_up__19 = one_hot_sel_158396[0] & nor_158451;
  assign exp__41 = exp__40 & sign_ext_157977;
  assign do_round_up__42 = one_hot_sel_158402[0] & nor_158456;
  assign exp__93 = exp__91 & sign_ext_158460;
  assign x_fraction__161 = x_fraction__159 & {24{ne_158434}};
  assign result_sign__804 = 1'h0;
  assign result_sign__805 = 1'h0;
  assign do_round_up__81 = one_hot_sel_158411[0] & nor_158464;
  assign exp__175 = exp__173 & sign_ext_157985;
  assign do_round_up__120 = one_hot_sel_158417[0] & nor_158469;
  assign exp__257 = exp__255 & sign_ext_158473;
  assign x_fraction__449 = x_fraction__447 & {24{ne_158447}};
  assign result_sign__806 = 1'h0;
  assign result_sign__807 = 1'h0;
  assign sel_158502 = do_round_up__19 ? {add_158453, nor_158451} : {result_sign__1116, one_hot_sel_158396, nor_158451};
  assign sel_158504 = do_round_up__42 ? {add_158458, nor_158456} : {result_sign__1117, one_hot_sel_158402, nor_158456};
  assign concat_158506 = {x_fraction__161, result_sign__804};
  assign concat_158507 = {result_sign__805, x_fraction__161};
  assign sel_158508 = do_round_up__81 ? {add_158466, nor_158464} : {result_sign__1118, one_hot_sel_158411, nor_158464};
  assign sel_158510 = do_round_up__120 ? {add_158471, nor_158469} : {result_sign__1119, one_hot_sel_158417, nor_158469};
  assign concat_158512 = {x_fraction__449, result_sign__806};
  assign concat_158513 = {result_sign__807, x_fraction__449};
  assign result_sign__391 = 1'h0;
  assign x_bexp__648 = 8'h00;
  assign rounding_carry__9 = sel_158502[25];
  assign sel_158517 = $signed(exp__41) <= $signed(10'h000) ? concat_158013 : concat_158012;
  assign result_sign__486 = 1'h0;
  assign x_bexp__649 = 8'h00;
  assign rounding_carry__20 = sel_158504[25];
  assign sel_158521 = $signed(exp__93) <= $signed(10'h000) ? concat_158507 : concat_158506;
  assign result_sign__581 = 1'h0;
  assign x_bexp__650 = 8'h00;
  assign rounding_carry__39 = sel_158508[25];
  assign sel_158525 = $signed(exp__175) <= $signed(10'h000) ? concat_158019 : concat_158018;
  assign result_sign__685 = 1'h0;
  assign x_bexp__651 = 8'h00;
  assign rounding_carry__58 = sel_158510[25];
  assign sel_158529 = $signed(exp__257) <= $signed(10'h000) ? concat_158513 : concat_158512;
  assign result_sign__929 = 1'h0;
  assign fraction__95 = sel_158517[23:1];
  assign result_sign__935 = 1'h0;
  assign fraction__208 = sel_158521[23:1];
  assign result_sign__941 = 1'h0;
  assign fraction__387 = sel_158525[23:1];
  assign result_sign__949 = 1'h0;
  assign fraction__566 = sel_158529[23:1];
  assign result_sign__392 = 1'h0;
  assign add_158547 = {result_sign__391, result_exp__29} + {x_bexp__648, rounding_carry__9};
  assign fraction__96 = {result_sign__929, fraction__95};
  assign result_sign__487 = 1'h0;
  assign add_158553 = {result_sign__486, result_exp__65} + {x_bexp__649, rounding_carry__20};
  assign fraction__210 = {result_sign__935, fraction__208};
  assign result_sign__582 = 1'h0;
  assign add_158559 = {result_sign__581, result_exp__125} + {x_bexp__650, rounding_carry__39};
  assign fraction__389 = {result_sign__941, fraction__387};
  assign result_sign__686 = 1'h0;
  assign add_158565 = {result_sign__685, result_exp__185} + {x_bexp__651, rounding_carry__58};
  assign fraction__568 = {result_sign__949, fraction__566};
  assign do_round_up__20 = sel_158517[0] & sel_158517[1];
  assign add_158576 = fraction__96 + 24'h00_0001;
  assign do_round_up__44 = sel_158521[0] & sel_158521[1];
  assign add_158583 = fraction__210 + 24'h00_0001;
  assign do_round_up__83 = sel_158525[0] & sel_158525[1];
  assign add_158590 = fraction__389 + 24'h00_0001;
  assign do_round_up__122 = sel_158529[0] & sel_158529[1];
  assign add_158597 = fraction__568 + 24'h00_0001;
  assign add_158598 = {result_sign__392, add_158547} + 10'h001;
  assign fraction__97 = do_round_up__20 ? add_158576 : fraction__96;
  assign add_158603 = {result_sign__487, add_158553} + 10'h001;
  assign fraction__212 = do_round_up__44 ? add_158583 : fraction__210;
  assign add_158608 = {result_sign__582, add_158559} + 10'h001;
  assign fraction__391 = do_round_up__83 ? add_158590 : fraction__389;
  assign add_158613 = {result_sign__686, add_158565} + 10'h001;
  assign fraction__570 = do_round_up__122 ? add_158597 : fraction__568;
  assign wide_exponent__27 = add_158598 - {5'h00, encode_158292};
  assign add_158621 = exp__41 + 10'h001;
  assign wide_exponent__58 = add_158603 - {5'h00, encode_158293};
  assign add_158625 = exp__93 + 10'h001;
  assign wide_exponent__115 = add_158608 - {5'h00, encode_158294};
  assign add_158629 = exp__175 + 10'h001;
  assign wide_exponent__172 = add_158613 - {5'h00, encode_158295};
  assign add_158633 = exp__257 + 10'h001;
  assign wide_exponent__28 = wide_exponent__27 & {10{fraction__89[28:3] != 26'h000_0000}};
  assign exp__43 = fraction__97[23] ? add_158621 : exp__41;
  assign wide_exponent__60 = wide_exponent__58 & {10{fraction__196[28:3] != 26'h000_0000}};
  assign exp__97 = fraction__212[23] ? add_158625 : exp__93;
  assign wide_exponent__117 = wide_exponent__115 & {10{fraction__375[28:3] != 26'h000_0000}};
  assign exp__179 = fraction__391[23] ? add_158629 : exp__175;
  assign wide_exponent__174 = wide_exponent__172 & {10{fraction__554[28:3] != 26'h000_0000}};
  assign exp__261 = fraction__570[23] ? add_158633 : exp__257;
  assign result_exp__30 = exp__43[8:0];
  assign result_exp__67 = exp__97[8:0];
  assign result_exp__127 = exp__179[8:0];
  assign result_exp__187 = exp__261[8:0];
  assign result_exp__31 = result_exp__30 & {9{$signed(exp__43) > $signed(10'h000)}};
  assign high_exp__146 = 8'hff;
  assign result_fraction__548 = 23'h00_0000;
  assign result_fraction__547 = 23'h00_0000;
  assign result_exp__69 = result_exp__67 & {9{$signed(exp__97) > $signed(10'h000)}};
  assign result_exp__129 = result_exp__127 & {9{$signed(exp__179) > $signed(10'h000)}};
  assign high_exp__280 = 8'hff;
  assign result_fraction__682 = 23'h00_0000;
  assign result_fraction__681 = 23'h00_0000;
  assign result_exp__189 = result_exp__187 & {9{$signed(exp__261) > $signed(10'h000)}};
  assign wide_exponent__29 = wide_exponent__28[8:0] & {9{~wide_exponent__28[9]}};
  assign result_fraction__770 = 23'h00_0000;
  assign result_fraction__483 = 23'h00_0000;
  assign wide_exponent__62 = wide_exponent__60[8:0] & {9{~wide_exponent__60[9]}};
  assign result_fraction__803 = 23'h00_0000;
  assign result_fraction__546 = 23'h00_0000;
  assign is_result_nan__45 = x_bexp__157 == high_exp__146;
  assign ne_158692 = x_fraction__157 != result_fraction__548;
  assign wide_exponent__119 = wide_exponent__117[8:0] & {9{~wide_exponent__117[9]}};
  assign result_fraction__836 = 23'h00_0000;
  assign result_fraction__613 = 23'h00_0000;
  assign wide_exponent__176 = wide_exponent__174[8:0] & {9{~wide_exponent__174[9]}};
  assign result_fraction__869 = 23'h00_0000;
  assign result_fraction__680 = 23'h00_0000;
  assign is_result_nan__123 = x_bexp__445 == high_exp__280;
  assign ne_158703 = x_fraction__445 != result_fraction__682;
  assign ne_158707 = result_fraction__56 != result_fraction__770;
  assign and_reduce_158711 = &result_exp__31[7:0];
  assign ne_158713 = result_fraction__122 != result_fraction__803;
  assign is_result_nan__44 = is_result_nan__45 & ne_158692;
  assign has_inf_arg__24 = is_result_nan__45 & x_fraction__157 == result_fraction__547;
  assign and_reduce_158719 = &result_exp__69[7:0];
  assign ne_158721 = result_fraction__239 != result_fraction__836;
  assign and_reduce_158725 = &result_exp__129[7:0];
  assign ne_158727 = result_fraction__356 != result_fraction__869;
  assign is_result_nan__122 = is_result_nan__123 & ne_158703;
  assign has_inf_arg__64 = is_result_nan__123 & x_fraction__445 == result_fraction__681;
  assign and_reduce_158733 = &result_exp__189[7:0];
  assign is_result_nan__19 = or_158158 & ne_158707;
  assign is_operand_inf__9 = or_158158 & result_fraction__56 == result_fraction__483;
  assign and_reduce_158740 = &wide_exponent__29[7:0];
  assign high_exp__83 = 8'hff;
  assign is_result_nan__42 = or_158162 & ne_158713;
  assign is_operand_inf__20 = or_158162 & result_fraction__122 == result_fraction__546;
  assign and_reduce_158749 = &wide_exponent__62[7:0];
  assign high_exp__147 = 8'hff;
  assign is_result_nan__81 = or_158166 & ne_158721;
  assign is_operand_inf__39 = or_158166 & result_fraction__239 == result_fraction__613;
  assign and_reduce_158758 = &wide_exponent__119[7:0];
  assign high_exp__212 = 8'hff;
  assign is_result_nan__120 = or_158170 & ne_158727;
  assign is_operand_inf__58 = or_158170 & result_fraction__356 == result_fraction__680;
  assign and_reduce_158767 = &wide_exponent__176[7:0];
  assign high_exp__281 = 8'hff;
  assign fraction_shift__29 = 3'h3;
  assign fraction_shift__28 = 3'h4;
  assign is_subnormal__10 = $signed(exp__43) <= $signed(10'h000);
  assign high_exp__82 = 8'hff;
  assign result_exp__32 = is_result_nan__40 | has_inf_arg__21 | result_exp__31[8] | and_reduce_158711 ? high_exp__83 : result_exp__31[7:0];
  assign fraction_shift__385 = 3'h3;
  assign fraction_shift__263 = 3'h4;
  assign is_subnormal__23 = $signed(exp__97) <= $signed(10'h000);
  assign high_exp__145 = 8'hff;
  assign result_exp__71 = is_result_nan__44 | has_inf_arg__24 | result_exp__69[8] | and_reduce_158719 ? high_exp__147 : result_exp__69[7:0];
  assign fraction_shift__403 = 3'h3;
  assign fraction_shift__298 = 3'h4;
  assign is_subnormal__43 = $signed(exp__179) <= $signed(10'h000);
  assign high_exp__211 = 8'hff;
  assign result_exp__131 = is_result_nan__118 | has_inf_arg__61 | result_exp__129[8] | and_reduce_158725 ? high_exp__212 : result_exp__129[7:0];
  assign fraction_shift__421 = 3'h3;
  assign fraction_shift__333 = 3'h4;
  assign is_subnormal__63 = $signed(exp__261) <= $signed(10'h000);
  assign high_exp__279 = 8'hff;
  assign result_exp__191 = is_result_nan__122 | has_inf_arg__64 | result_exp__189[8] | and_reduce_158733 ? high_exp__281 : result_exp__189[7:0];
  assign result_exp__6 = {8{is_result_nan__3}};
  assign rounded_fraction__9 = {sel_158502, 2'h0};
  assign fraction_shift__30 = rounding_carry__9 ? fraction_shift__28 : fraction_shift__29;
  assign result_sign__393 = 1'h0;
  assign result_exponent__10 = is_result_nan__19 | is_operand_inf__9 | wide_exponent__29[8] | and_reduce_158740 ? high_exp__82 : wide_exponent__29[7:0];
  assign result_sign__394 = 1'h0;
  assign result_exp__72 = {8{is_result_nan__45}};
  assign rounded_fraction__20 = {sel_158504, 2'h0};
  assign fraction_shift__62 = rounding_carry__20 ? fraction_shift__263 : fraction_shift__385;
  assign result_sign__488 = 1'h0;
  assign result_exponent__20 = is_result_nan__42 | is_operand_inf__20 | wide_exponent__62[8] | and_reduce_158749 ? high_exp__145 : wide_exponent__62[7:0];
  assign result_sign__489 = 1'h0;
  assign result_exp__132 = {8{is_result_nan__84}};
  assign rounded_fraction__39 = {sel_158508, 2'h0};
  assign fraction_shift__119 = rounding_carry__39 ? fraction_shift__298 : fraction_shift__403;
  assign result_sign__583 = 1'h0;
  assign result_exponent__39 = is_result_nan__81 | is_operand_inf__39 | wide_exponent__119[8] | and_reduce_158758 ? high_exp__211 : wide_exponent__119[7:0];
  assign result_sign__584 = 1'h0;
  assign result_exp__192 = {8{is_result_nan__123}};
  assign rounded_fraction__58 = {sel_158510, 2'h0};
  assign fraction_shift__176 = rounding_carry__58 ? fraction_shift__333 : fraction_shift__421;
  assign result_sign__687 = 1'h0;
  assign result_exponent__58 = is_result_nan__120 | is_operand_inf__58 | wide_exponent__176[8] | and_reduce_158767 ? high_exp__279 : wide_exponent__176[7:0];
  assign result_sign__688 = 1'h0;
  assign result_sign__395 = 1'h0;
  assign shrl_158840 = rounded_fraction__9 >> fraction_shift__30;
  assign concat_158843 = {result_sign__393, result_exponent__10};
  assign result_sign__490 = 1'h0;
  assign shrl_158847 = rounded_fraction__20 >> fraction_shift__62;
  assign concat_158850 = {result_sign__488, result_exponent__20};
  assign result_sign__585 = 1'h0;
  assign shrl_158854 = rounded_fraction__39 >> fraction_shift__119;
  assign concat_158857 = {result_sign__583, result_exponent__39};
  assign concat_158858 = {result_sign__584, ~result_exp__131};
  assign result_sign__689 = 1'h0;
  assign shrl_158861 = rounded_fraction__58 >> fraction_shift__176;
  assign concat_158864 = {result_sign__687, result_exponent__58};
  assign concat_158865 = {result_sign__688, ~result_exp__191};
  assign result_fraction__57 = shrl_158840[22:0];
  assign result_fraction__60 = fraction__97[22:0];
  assign sum__10 = concat_158843 + {result_sign__394, ~result_exp__32};
  assign result_fraction__124 = shrl_158847[22:0];
  assign result_fraction__130 = fraction__212[22:0];
  assign sum__22 = concat_158850 + {result_sign__489, ~result_exp__71};
  assign concat_158878 = {result_sign__585, ~result_exp__132};
  assign result_fraction__241 = shrl_158854[22:0];
  assign result_fraction__247 = fraction__391[22:0];
  assign sum__41 = concat_158857 + concat_158858;
  assign concat_158884 = {result_sign__689, ~result_exp__192};
  assign result_fraction__358 = shrl_158861[22:0];
  assign result_fraction__364 = fraction__570[22:0];
  assign sum__60 = concat_158864 + concat_158865;
  assign sum__2 = concat_158843 + {result_sign__395, ~result_exp__6};
  assign result_fraction__58 = result_fraction__57 & {23{~(is_operand_inf__9 | wide_exponent__29[8] | and_reduce_158740 | ~((|wide_exponent__29[8:1]) | wide_exponent__29[0]))}};
  assign nan_fraction__81 = 23'h40_0000;
  assign result_fraction__61 = result_fraction__60 & {23{~(has_inf_arg__21 | result_exp__31[8] | and_reduce_158711 | is_subnormal__10)}};
  assign nan_fraction__82 = 23'h40_0000;
  assign sum__23 = concat_158850 + {result_sign__490, ~result_exp__72};
  assign result_fraction__126 = result_fraction__124 & {23{~(is_operand_inf__20 | wide_exponent__62[8] | and_reduce_158749 | ~((|wide_exponent__62[8:1]) | wide_exponent__62[0]))}};
  assign nan_fraction__108 = 23'h40_0000;
  assign result_fraction__132 = result_fraction__130 & {23{~(has_inf_arg__24 | result_exp__69[8] | and_reduce_158719 | is_subnormal__23)}};
  assign nan_fraction__109 = 23'h40_0000;
  assign sum__42 = concat_158857 + concat_158878;
  assign result_fraction__243 = result_fraction__241 & {23{~(is_operand_inf__39 | wide_exponent__119[8] | and_reduce_158758 | ~((|wide_exponent__119[8:1]) | wide_exponent__119[0]))}};
  assign nan_fraction__135 = 23'h40_0000;
  assign result_fraction__249 = result_fraction__247 & {23{~(has_inf_arg__61 | result_exp__129[8] | and_reduce_158725 | is_subnormal__43)}};
  assign nan_fraction__136 = 23'h40_0000;
  assign sum__61 = concat_158864 + concat_158884;
  assign result_fraction__360 = result_fraction__358 & {23{~(is_operand_inf__58 | wide_exponent__176[8] | and_reduce_158767 | ~((|wide_exponent__176[8:1]) | wide_exponent__176[0]))}};
  assign nan_fraction__164 = 23'h40_0000;
  assign result_fraction__366 = result_fraction__364 & {23{~(has_inf_arg__64 | result_exp__189[8] | and_reduce_158733 | is_subnormal__63)}};
  assign nan_fraction__165 = 23'h40_0000;
  assign result_fraction__59 = is_result_nan__19 ? nan_fraction__81 : result_fraction__58;
  assign result_fraction__62 = is_result_nan__40 ? nan_fraction__82 : result_fraction__61;
  assign prod_bexp__42 = sum__10[8] ? result_exp__32 : result_exponent__10;
  assign x_bexp__674 = 8'h00;
  assign result_fraction__128 = is_result_nan__42 ? nan_fraction__108 : result_fraction__126;
  assign result_fraction__134 = is_result_nan__44 ? nan_fraction__109 : result_fraction__132;
  assign prod_bexp__83 = sum__22[8] ? result_exp__71 : result_exponent__20;
  assign x_bexp__675 = 8'h00;
  assign result_fraction__245 = is_result_nan__81 ? nan_fraction__135 : result_fraction__243;
  assign result_fraction__251 = is_result_nan__118 ? nan_fraction__136 : result_fraction__249;
  assign prod_bexp__155 = sum__41[8] ? result_exp__131 : result_exponent__39;
  assign x_bexp__676 = 8'h00;
  assign result_fraction__362 = is_result_nan__120 ? nan_fraction__164 : result_fraction__360;
  assign result_fraction__368 = is_result_nan__122 ? nan_fraction__165 : result_fraction__366;
  assign prod_bexp__227 = sum__60[8] ? result_exp__191 : result_exponent__58;
  assign x_bexp__677 = 8'h00;
  assign result_fraction__469 = {is_result_nan__3, 22'h00_0000};
  assign prod_bexp__6 = sum__2[8] ? result_exp__6 : result_exponent__10;
  assign x_bexp__678 = 8'h00;
  assign prod_fraction__30 = sum__10[8] ? result_fraction__62 : result_fraction__59;
  assign incremented_sum__78 = sum__10[7:0] + 8'h01;
  assign result_fraction__470 = {is_result_nan__45, 22'h00_0000};
  assign prod_bexp__84 = sum__23[8] ? result_exp__72 : result_exponent__20;
  assign x_bexp__679 = 8'h00;
  assign prod_fraction__61 = sum__22[8] ? result_fraction__134 : result_fraction__128;
  assign incremented_sum__96 = sum__22[7:0] + 8'h01;
  assign result_fraction__471 = {is_result_nan__84, 22'h00_0000};
  assign prod_bexp__156 = sum__42[8] ? result_exp__132 : result_exponent__39;
  assign x_bexp__680 = 8'h00;
  assign prod_fraction__115 = sum__41[8] ? result_fraction__251 : result_fraction__245;
  assign incremented_sum__114 = sum__41[7:0] + 8'h01;
  assign result_fraction__472 = {is_result_nan__123, 22'h00_0000};
  assign prod_bexp__228 = sum__61[8] ? result_exp__192 : result_exponent__58;
  assign x_bexp__681 = 8'h00;
  assign prod_fraction__169 = sum__60[8] ? result_fraction__368 : result_fraction__362;
  assign incremented_sum__132 = sum__60[7:0] + 8'h01;
  assign prod_fraction__4 = sum__2[8] ? result_fraction__469 : result_fraction__59;
  assign incremented_sum__79 = sum__2[7:0] + 8'h01;
  assign wide_y__20 = {2'h1, prod_fraction__30, 3'h0};
  assign x_bexpbs_difference__11 = sum__10[8] ? incremented_sum__78 : ~sum__10[7:0];
  assign prod_fraction__62 = sum__23[8] ? result_fraction__470 : result_fraction__128;
  assign incremented_sum__97 = sum__23[7:0] + 8'h01;
  assign wide_y__43 = {2'h1, prod_fraction__61, 3'h0};
  assign x_bexpbs_difference__21 = sum__22[8] ? incremented_sum__96 : ~sum__22[7:0];
  assign prod_fraction__116 = sum__42[8] ? result_fraction__471 : result_fraction__245;
  assign incremented_sum__115 = sum__42[7:0] + 8'h01;
  assign wide_y__81 = {2'h1, prod_fraction__115, 3'h0};
  assign x_bexpbs_difference__39 = sum__41[8] ? incremented_sum__114 : ~sum__41[7:0];
  assign prod_fraction__170 = sum__61[8] ? result_fraction__472 : result_fraction__362;
  assign incremented_sum__133 = sum__61[7:0] + 8'h01;
  assign wide_y__119 = {2'h1, prod_fraction__169, 3'h0};
  assign x_bexpbs_difference__57 = sum__60[8] ? incremented_sum__132 : ~sum__60[7:0];
  assign wide_y__3 = {2'h1, prod_fraction__4, 3'h0};
  assign x_bexpbs_difference__2 = sum__2[8] ? incremented_sum__79 : ~sum__2[7:0];
  assign has_pos_inf__9 = ~(ne_158707 | result_sign__46);
  assign x_bexp__86 = sum__10[8] ? result_exponent__10 : result_exp__32;
  assign x_bexp__682 = 8'h00;
  assign wide_y__21 = wide_y__20 & {28{prod_bexp__42 != x_bexp__674}};
  assign sub_159038 = 8'h1c - x_bexpbs_difference__11;
  assign wide_y__44 = {2'h1, prod_fraction__62, 3'h0};
  assign x_bexpbs_difference__22 = sum__23[8] ? incremented_sum__97 : ~sum__23[7:0];
  assign has_pos_inf__20 = ~(ne_158713 | result_sign__100);
  assign x_bexp__171 = sum__22[8] ? result_exponent__20 : result_exp__71;
  assign x_bexp__683 = 8'h00;
  assign wide_y__45 = wide_y__43 & {28{prod_bexp__83 != x_bexp__675}};
  assign sub_159047 = 8'h1c - x_bexpbs_difference__21;
  assign wide_y__82 = {2'h1, prod_fraction__116, 3'h0};
  assign x_bexpbs_difference__40 = sum__42[8] ? incremented_sum__115 : ~sum__42[7:0];
  assign has_pos_inf__39 = ~(ne_158721 | result_sign__197);
  assign x_bexp__315 = sum__41[8] ? result_exponent__39 : result_exp__131;
  assign x_bexp__684 = 8'h00;
  assign wide_y__83 = wide_y__81 & {28{prod_bexp__155 != x_bexp__676}};
  assign sub_159056 = 8'h1c - x_bexpbs_difference__39;
  assign wide_y__120 = {2'h1, prod_fraction__170, 3'h0};
  assign x_bexpbs_difference__58 = sum__61[8] ? incremented_sum__133 : ~sum__61[7:0];
  assign has_pos_inf__58 = ~(ne_158727 | result_sign__294);
  assign x_bexp__459 = sum__60[8] ? result_exponent__58 : result_exp__191;
  assign x_bexp__685 = 8'h00;
  assign wide_y__121 = wide_y__119 & {28{prod_bexp__227 != x_bexp__677}};
  assign sub_159065 = 8'h1c - x_bexpbs_difference__57;
  assign x_bexp__14 = sum__2[8] ? result_exponent__10 : result_exp__6;
  assign x_bexp__686 = 8'h00;
  assign wide_y__4 = wide_y__3 & {28{prod_bexp__6 != x_bexp__678}};
  assign sub_159069 = 8'h1c - x_bexpbs_difference__2;
  assign x_fraction__86 = sum__10[8] ? result_fraction__59 : result_fraction__62;
  assign dropped__10 = sub_159038 >= 8'h1c ? 28'h000_0000 : wide_y__21 << sub_159038;
  assign x_bexp__172 = sum__23[8] ? result_exponent__20 : result_exp__72;
  assign x_bexp__687 = 8'h00;
  assign wide_y__46 = wide_y__44 & {28{prod_bexp__84 != x_bexp__679}};
  assign sub_159079 = 8'h1c - x_bexpbs_difference__22;
  assign x_sign__41 = array_index_158318[31:31];
  assign x_fraction__171 = sum__22[8] ? result_fraction__128 : result_fraction__134;
  assign dropped__22 = sub_159047 >= 8'h1c ? 28'h000_0000 : wide_y__45 << sub_159047;
  assign x_bexp__316 = sum__42[8] ? result_exponent__39 : result_exp__132;
  assign x_bexp__688 = 8'h00;
  assign wide_y__84 = wide_y__82 & {28{prod_bexp__156 != x_bexp__680}};
  assign sub_159090 = 8'h1c - x_bexpbs_difference__40;
  assign x_fraction__315 = sum__41[8] ? result_fraction__245 : result_fraction__251;
  assign dropped__41 = sub_159056 >= 8'h1c ? 28'h000_0000 : wide_y__83 << sub_159056;
  assign x_bexp__460 = sum__61[8] ? result_exponent__58 : result_exp__192;
  assign x_bexp__689 = 8'h00;
  assign wide_y__122 = wide_y__120 & {28{prod_bexp__228 != x_bexp__681}};
  assign sub_159100 = 8'h1c - x_bexpbs_difference__58;
  assign x_sign__113 = array_index_158331[31:31];
  assign x_fraction__459 = sum__60[8] ? result_fraction__362 : result_fraction__368;
  assign dropped__60 = sub_159065 >= 8'h1c ? 28'h000_0000 : wide_y__121 << sub_159065;
  assign high_exp__479 = 8'hff;
  assign x_fraction__14 = sum__2[8] ? result_fraction__59 : result_fraction__469;
  assign dropped__2 = sub_159069 >= 8'h1c ? 28'h000_0000 : wide_y__4 << sub_159069;
  assign result_sign__48 = is_operand_inf__9 ? ~has_pos_inf__9 : result_sign__47;
  assign wide_x__20 = {2'h1, x_fraction__86, 3'h0};
  assign high_exp__481 = 8'hff;
  assign x_fraction__172 = sum__23[8] ? result_fraction__128 : result_fraction__470;
  assign dropped__23 = sub_159079 >= 8'h1c ? 28'h000_0000 : wide_y__46 << sub_159079;
  assign nand_159126 = ~(is_result_nan__45 & ne_158692);
  assign result_sign__108 = ~x_sign__41;
  assign result_sign__104 = is_operand_inf__20 ? ~has_pos_inf__20 : result_sign__102;
  assign wide_x__43 = {2'h1, x_fraction__171, 3'h0};
  assign high_exp__483 = 8'hff;
  assign x_fraction__316 = sum__42[8] ? result_fraction__245 : result_fraction__471;
  assign dropped__42 = sub_159090 >= 8'h1c ? 28'h000_0000 : wide_y__84 << sub_159090;
  assign result_sign__201 = is_operand_inf__39 ? ~has_pos_inf__39 : result_sign__199;
  assign wide_x__81 = {2'h1, x_fraction__315, 3'h0};
  assign high_exp__486 = 8'hff;
  assign x_fraction__460 = sum__61[8] ? result_fraction__362 : result_fraction__472;
  assign dropped__61 = sub_159100 >= 8'h1c ? 28'h000_0000 : wide_y__122 << sub_159100;
  assign nand_159152 = ~(is_result_nan__123 & ne_158703);
  assign result_sign__302 = ~x_sign__113;
  assign result_sign__298 = is_operand_inf__58 ? ~has_pos_inf__58 : result_sign__296;
  assign wide_x__119 = {2'h1, x_fraction__459, 3'h0};
  assign wide_x__3 = {2'h1, x_fraction__14, 3'h0};
  assign result_sign__49 = ~(or_158158 & ne_158707) & result_sign__48;
  assign wide_x__21 = wide_x__20 & {28{x_bexp__86 != x_bexp__682}};
  assign wide_x__44 = {2'h1, x_fraction__172, 3'h0};
  assign result_sign__110 = nand_159126 & result_sign__108;
  assign result_sign__106 = ~(or_158162 & ne_158713) & result_sign__104;
  assign wide_x__45 = wide_x__43 & {28{x_bexp__171 != x_bexp__683}};
  assign wide_x__82 = {2'h1, x_fraction__316, 3'h0};
  assign result_sign__203 = ~(or_158166 & ne_158721) & result_sign__201;
  assign wide_x__83 = wide_x__81 & {28{x_bexp__315 != x_bexp__684}};
  assign wide_x__120 = {2'h1, x_fraction__460, 3'h0};
  assign result_sign__304 = nand_159152 & result_sign__302;
  assign result_sign__300 = ~(or_158170 & ne_158727) & result_sign__298;
  assign wide_x__121 = wide_x__119 & {28{x_bexp__459 != x_bexp__685}};
  assign result_sign__7 = x_bexp__145 != high_exp__479 & x_sign__37;
  assign wide_x__4 = wide_x__3 & {28{x_bexp__14 != x_bexp__686}};
  assign x_sign__22 = sum__10[8] ? result_sign__49 : result_sign__100;
  assign prod_sign__10 = sum__10[8] ? result_sign__100 : result_sign__49;
  assign neg_159204 = -wide_x__21;
  assign sticky__32 = {27'h000_0000, dropped__10[27:3] != 25'h000_0000};
  assign result_sign__111 = x_bexp__157 != high_exp__481 & x_sign__41;
  assign wide_x__46 = wide_x__44 & {28{x_bexp__172 != x_bexp__687}};
  assign x_sign__43 = sum__22[8] ? result_sign__106 : result_sign__110;
  assign prod_sign__21 = sum__22[8] ? result_sign__110 : result_sign__106;
  assign neg_159213 = -wide_x__45;
  assign sticky__70 = {27'h000_0000, dropped__22[27:3] != 25'h000_0000};
  assign result_sign__208 = x_bexp__433 != high_exp__483 & x_sign__109;
  assign wide_x__84 = wide_x__82 & {28{x_bexp__316 != x_bexp__688}};
  assign x_sign__79 = sum__41[8] ? result_sign__203 : result_sign__294;
  assign prod_sign__39 = sum__41[8] ? result_sign__294 : result_sign__203;
  assign neg_159222 = -wide_x__83;
  assign sticky__129 = {27'h000_0000, dropped__41[27:3] != 25'h000_0000};
  assign result_sign__305 = x_bexp__445 != high_exp__486 & x_sign__113;
  assign wide_x__122 = wide_x__120 & {28{x_bexp__460 != x_bexp__689}};
  assign x_sign__115 = sum__60[8] ? result_sign__300 : result_sign__304;
  assign prod_sign__57 = sum__60[8] ? result_sign__304 : result_sign__300;
  assign neg_159231 = -wide_x__121;
  assign sticky__188 = {27'h000_0000, dropped__60[27:3] != 25'h000_0000};
  assign x_sign__4 = sum__2[8] ? result_sign__49 : result_sign__7;
  assign prod_sign__2 = sum__2[8] ? result_sign__7 : result_sign__49;
  assign neg_159236 = -wide_x__4;
  assign sticky__6 = {27'h000_0000, dropped__2[27:3] != 25'h000_0000};
  assign xddend_y__10 = (x_bexpbs_difference__11 >= 8'h1c ? 28'h000_0000 : wide_y__21 >> x_bexpbs_difference__11) | sticky__32;
  assign x_sign__44 = sum__23[8] ? result_sign__106 : result_sign__111;
  assign prod_sign__22 = sum__23[8] ? result_sign__111 : result_sign__106;
  assign neg_159245 = -wide_x__46;
  assign sticky__71 = {27'h000_0000, dropped__23[27:3] != 25'h000_0000};
  assign xddend_y__21 = (x_bexpbs_difference__21 >= 8'h1c ? 28'h000_0000 : wide_y__45 >> x_bexpbs_difference__21) | sticky__70;
  assign x_sign__80 = sum__42[8] ? result_sign__203 : result_sign__208;
  assign prod_sign__40 = sum__42[8] ? result_sign__208 : result_sign__203;
  assign neg_159254 = -wide_x__84;
  assign sticky__130 = {27'h000_0000, dropped__42[27:3] != 25'h000_0000};
  assign xddend_y__39 = (x_bexpbs_difference__39 >= 8'h1c ? 28'h000_0000 : wide_y__83 >> x_bexpbs_difference__39) | sticky__129;
  assign x_sign__116 = sum__61[8] ? result_sign__300 : result_sign__305;
  assign prod_sign__58 = sum__61[8] ? result_sign__305 : result_sign__300;
  assign neg_159263 = -wide_x__122;
  assign sticky__189 = {27'h000_0000, dropped__61[27:3] != 25'h000_0000};
  assign xddend_y__57 = (x_bexpbs_difference__57 >= 8'h1c ? 28'h000_0000 : wide_y__121 >> x_bexpbs_difference__57) | sticky__188;
  assign xddend_y__2 = (x_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : wide_y__4 >> x_bexpbs_difference__2) | sticky__6;
  assign sel_159274 = x_sign__22 ^ prod_sign__10 ? neg_159204[27:3] : wide_x__21[27:3];
  assign result_sign__964 = 1'h0;
  assign xddend_y__22 = (x_bexpbs_difference__22 >= 8'h1c ? 28'h000_0000 : wide_y__46 >> x_bexpbs_difference__22) | sticky__71;
  assign sel_159281 = x_sign__43 ^ prod_sign__21 ? neg_159213[27:3] : wide_x__45[27:3];
  assign result_sign__965 = 1'h0;
  assign xddend_y__40 = (x_bexpbs_difference__40 >= 8'h1c ? 28'h000_0000 : wide_y__84 >> x_bexpbs_difference__40) | sticky__130;
  assign sel_159288 = x_sign__79 ^ prod_sign__39 ? neg_159222[27:3] : wide_x__83[27:3];
  assign result_sign__966 = 1'h0;
  assign xddend_y__58 = (x_bexpbs_difference__58 >= 8'h1c ? 28'h000_0000 : wide_y__122 >> x_bexpbs_difference__58) | sticky__189;
  assign sel_159295 = x_sign__115 ^ prod_sign__57 ? neg_159231[27:3] : wide_x__121[27:3];
  assign result_sign__967 = 1'h0;
  assign sel_159298 = x_sign__4 ^ prod_sign__2 ? neg_159236[27:3] : wide_x__4[27:3];
  assign result_sign__968 = 1'h0;
  assign sel_159303 = x_sign__44 ^ prod_sign__22 ? neg_159245[27:3] : wide_x__46[27:3];
  assign result_sign__969 = 1'h0;
  assign sel_159308 = x_sign__80 ^ prod_sign__40 ? neg_159254[27:3] : wide_x__84[27:3];
  assign result_sign__970 = 1'h0;
  assign sel_159313 = x_sign__116 ^ prod_sign__58 ? neg_159263[27:3] : wide_x__122[27:3];
  assign result_sign__971 = 1'h0;
  assign add_159320 = {{1{sel_159274[24]}}, sel_159274} + {result_sign__964, xddend_y__10[27:3]};
  assign add_159323 = {{1{sel_159281[24]}}, sel_159281} + {result_sign__965, xddend_y__21[27:3]};
  assign add_159326 = {{1{sel_159288[24]}}, sel_159288} + {result_sign__966, xddend_y__39[27:3]};
  assign add_159329 = {{1{sel_159295[24]}}, sel_159295} + {result_sign__967, xddend_y__57[27:3]};
  assign add_159330 = {{1{sel_159298[24]}}, sel_159298} + {result_sign__968, xddend_y__2[27:3]};
  assign add_159333 = {{1{sel_159303[24]}}, sel_159303} + {result_sign__969, xddend_y__22[27:3]};
  assign add_159336 = {{1{sel_159308[24]}}, sel_159308} + {result_sign__970, xddend_y__40[27:3]};
  assign add_159339 = {{1{sel_159313[24]}}, sel_159313} + {result_sign__971, xddend_y__58[27:3]};
  assign concat_159344 = {add_159320[24:0], xddend_y__10[2:0]};
  assign concat_159347 = {add_159323[24:0], xddend_y__21[2:0]};
  assign concat_159350 = {add_159326[24:0], xddend_y__39[2:0]};
  assign concat_159353 = {add_159329[24:0], xddend_y__57[2:0]};
  assign concat_159354 = {add_159330[24:0], xddend_y__2[2:0]};
  assign concat_159357 = {add_159333[24:0], xddend_y__22[2:0]};
  assign concat_159360 = {add_159336[24:0], xddend_y__40[2:0]};
  assign concat_159363 = {add_159339[24:0], xddend_y__58[2:0]};
  assign xbs_fraction__10 = add_159320[25] ? -concat_159344 : concat_159344;
  assign xbs_fraction__21 = add_159323[25] ? -concat_159347 : concat_159347;
  assign xbs_fraction__39 = add_159326[25] ? -concat_159350 : concat_159350;
  assign xbs_fraction__57 = add_159329[25] ? -concat_159353 : concat_159353;
  assign xbs_fraction__2 = add_159330[25] ? -concat_159354 : concat_159354;
  assign reverse_159379 = {xbs_fraction__10[0], xbs_fraction__10[1], xbs_fraction__10[2], xbs_fraction__10[3], xbs_fraction__10[4], xbs_fraction__10[5], xbs_fraction__10[6], xbs_fraction__10[7], xbs_fraction__10[8], xbs_fraction__10[9], xbs_fraction__10[10], xbs_fraction__10[11], xbs_fraction__10[12], xbs_fraction__10[13], xbs_fraction__10[14], xbs_fraction__10[15], xbs_fraction__10[16], xbs_fraction__10[17], xbs_fraction__10[18], xbs_fraction__10[19], xbs_fraction__10[20], xbs_fraction__10[21], xbs_fraction__10[22], xbs_fraction__10[23], xbs_fraction__10[24], xbs_fraction__10[25], xbs_fraction__10[26], xbs_fraction__10[27]};
  assign xbs_fraction__22 = add_159333[25] ? -concat_159357 : concat_159357;
  assign reverse_159381 = {xbs_fraction__21[0], xbs_fraction__21[1], xbs_fraction__21[2], xbs_fraction__21[3], xbs_fraction__21[4], xbs_fraction__21[5], xbs_fraction__21[6], xbs_fraction__21[7], xbs_fraction__21[8], xbs_fraction__21[9], xbs_fraction__21[10], xbs_fraction__21[11], xbs_fraction__21[12], xbs_fraction__21[13], xbs_fraction__21[14], xbs_fraction__21[15], xbs_fraction__21[16], xbs_fraction__21[17], xbs_fraction__21[18], xbs_fraction__21[19], xbs_fraction__21[20], xbs_fraction__21[21], xbs_fraction__21[22], xbs_fraction__21[23], xbs_fraction__21[24], xbs_fraction__21[25], xbs_fraction__21[26], xbs_fraction__21[27]};
  assign xbs_fraction__40 = add_159336[25] ? -concat_159360 : concat_159360;
  assign reverse_159383 = {xbs_fraction__39[0], xbs_fraction__39[1], xbs_fraction__39[2], xbs_fraction__39[3], xbs_fraction__39[4], xbs_fraction__39[5], xbs_fraction__39[6], xbs_fraction__39[7], xbs_fraction__39[8], xbs_fraction__39[9], xbs_fraction__39[10], xbs_fraction__39[11], xbs_fraction__39[12], xbs_fraction__39[13], xbs_fraction__39[14], xbs_fraction__39[15], xbs_fraction__39[16], xbs_fraction__39[17], xbs_fraction__39[18], xbs_fraction__39[19], xbs_fraction__39[20], xbs_fraction__39[21], xbs_fraction__39[22], xbs_fraction__39[23], xbs_fraction__39[24], xbs_fraction__39[25], xbs_fraction__39[26], xbs_fraction__39[27]};
  assign xbs_fraction__58 = add_159339[25] ? -concat_159363 : concat_159363;
  assign reverse_159385 = {xbs_fraction__57[0], xbs_fraction__57[1], xbs_fraction__57[2], xbs_fraction__57[3], xbs_fraction__57[4], xbs_fraction__57[5], xbs_fraction__57[6], xbs_fraction__57[7], xbs_fraction__57[8], xbs_fraction__57[9], xbs_fraction__57[10], xbs_fraction__57[11], xbs_fraction__57[12], xbs_fraction__57[13], xbs_fraction__57[14], xbs_fraction__57[15], xbs_fraction__57[16], xbs_fraction__57[17], xbs_fraction__57[18], xbs_fraction__57[19], xbs_fraction__57[20], xbs_fraction__57[21], xbs_fraction__57[22], xbs_fraction__57[23], xbs_fraction__57[24], xbs_fraction__57[25], xbs_fraction__57[26], xbs_fraction__57[27]};
  assign reverse_159386 = {xbs_fraction__2[0], xbs_fraction__2[1], xbs_fraction__2[2], xbs_fraction__2[3], xbs_fraction__2[4], xbs_fraction__2[5], xbs_fraction__2[6], xbs_fraction__2[7], xbs_fraction__2[8], xbs_fraction__2[9], xbs_fraction__2[10], xbs_fraction__2[11], xbs_fraction__2[12], xbs_fraction__2[13], xbs_fraction__2[14], xbs_fraction__2[15], xbs_fraction__2[16], xbs_fraction__2[17], xbs_fraction__2[18], xbs_fraction__2[19], xbs_fraction__2[20], xbs_fraction__2[21], xbs_fraction__2[22], xbs_fraction__2[23], xbs_fraction__2[24], xbs_fraction__2[25], xbs_fraction__2[26], xbs_fraction__2[27]};
  assign one_hot_159387 = {reverse_159379[27:0] == 28'h000_0000, reverse_159379[27] && reverse_159379[26:0] == 27'h000_0000, reverse_159379[26] && reverse_159379[25:0] == 26'h000_0000, reverse_159379[25] && reverse_159379[24:0] == 25'h000_0000, reverse_159379[24] && reverse_159379[23:0] == 24'h00_0000, reverse_159379[23] && reverse_159379[22:0] == 23'h00_0000, reverse_159379[22] && reverse_159379[21:0] == 22'h00_0000, reverse_159379[21] && reverse_159379[20:0] == 21'h00_0000, reverse_159379[20] && reverse_159379[19:0] == 20'h0_0000, reverse_159379[19] && reverse_159379[18:0] == 19'h0_0000, reverse_159379[18] && reverse_159379[17:0] == 18'h0_0000, reverse_159379[17] && reverse_159379[16:0] == 17'h0_0000, reverse_159379[16] && reverse_159379[15:0] == 16'h0000, reverse_159379[15] && reverse_159379[14:0] == 15'h0000, reverse_159379[14] && reverse_159379[13:0] == 14'h0000, reverse_159379[13] && reverse_159379[12:0] == 13'h0000, reverse_159379[12] && reverse_159379[11:0] == 12'h000, reverse_159379[11] && reverse_159379[10:0] == 11'h000, reverse_159379[10] && reverse_159379[9:0] == 10'h000, reverse_159379[9] && reverse_159379[8:0] == 9'h000, reverse_159379[8] && reverse_159379[7:0] == 8'h00, reverse_159379[7] && reverse_159379[6:0] == 7'h00, reverse_159379[6] && reverse_159379[5:0] == 6'h00, reverse_159379[5] && reverse_159379[4:0] == 5'h00, reverse_159379[4] && reverse_159379[3:0] == 4'h0, reverse_159379[3] && reverse_159379[2:0] == 3'h0, reverse_159379[2] && reverse_159379[1:0] == 2'h0, reverse_159379[1] && !reverse_159379[0], reverse_159379[0]};
  assign reverse_159388 = {xbs_fraction__22[0], xbs_fraction__22[1], xbs_fraction__22[2], xbs_fraction__22[3], xbs_fraction__22[4], xbs_fraction__22[5], xbs_fraction__22[6], xbs_fraction__22[7], xbs_fraction__22[8], xbs_fraction__22[9], xbs_fraction__22[10], xbs_fraction__22[11], xbs_fraction__22[12], xbs_fraction__22[13], xbs_fraction__22[14], xbs_fraction__22[15], xbs_fraction__22[16], xbs_fraction__22[17], xbs_fraction__22[18], xbs_fraction__22[19], xbs_fraction__22[20], xbs_fraction__22[21], xbs_fraction__22[22], xbs_fraction__22[23], xbs_fraction__22[24], xbs_fraction__22[25], xbs_fraction__22[26], xbs_fraction__22[27]};
  assign one_hot_159389 = {reverse_159381[27:0] == 28'h000_0000, reverse_159381[27] && reverse_159381[26:0] == 27'h000_0000, reverse_159381[26] && reverse_159381[25:0] == 26'h000_0000, reverse_159381[25] && reverse_159381[24:0] == 25'h000_0000, reverse_159381[24] && reverse_159381[23:0] == 24'h00_0000, reverse_159381[23] && reverse_159381[22:0] == 23'h00_0000, reverse_159381[22] && reverse_159381[21:0] == 22'h00_0000, reverse_159381[21] && reverse_159381[20:0] == 21'h00_0000, reverse_159381[20] && reverse_159381[19:0] == 20'h0_0000, reverse_159381[19] && reverse_159381[18:0] == 19'h0_0000, reverse_159381[18] && reverse_159381[17:0] == 18'h0_0000, reverse_159381[17] && reverse_159381[16:0] == 17'h0_0000, reverse_159381[16] && reverse_159381[15:0] == 16'h0000, reverse_159381[15] && reverse_159381[14:0] == 15'h0000, reverse_159381[14] && reverse_159381[13:0] == 14'h0000, reverse_159381[13] && reverse_159381[12:0] == 13'h0000, reverse_159381[12] && reverse_159381[11:0] == 12'h000, reverse_159381[11] && reverse_159381[10:0] == 11'h000, reverse_159381[10] && reverse_159381[9:0] == 10'h000, reverse_159381[9] && reverse_159381[8:0] == 9'h000, reverse_159381[8] && reverse_159381[7:0] == 8'h00, reverse_159381[7] && reverse_159381[6:0] == 7'h00, reverse_159381[6] && reverse_159381[5:0] == 6'h00, reverse_159381[5] && reverse_159381[4:0] == 5'h00, reverse_159381[4] && reverse_159381[3:0] == 4'h0, reverse_159381[3] && reverse_159381[2:0] == 3'h0, reverse_159381[2] && reverse_159381[1:0] == 2'h0, reverse_159381[1] && !reverse_159381[0], reverse_159381[0]};
  assign reverse_159390 = {xbs_fraction__40[0], xbs_fraction__40[1], xbs_fraction__40[2], xbs_fraction__40[3], xbs_fraction__40[4], xbs_fraction__40[5], xbs_fraction__40[6], xbs_fraction__40[7], xbs_fraction__40[8], xbs_fraction__40[9], xbs_fraction__40[10], xbs_fraction__40[11], xbs_fraction__40[12], xbs_fraction__40[13], xbs_fraction__40[14], xbs_fraction__40[15], xbs_fraction__40[16], xbs_fraction__40[17], xbs_fraction__40[18], xbs_fraction__40[19], xbs_fraction__40[20], xbs_fraction__40[21], xbs_fraction__40[22], xbs_fraction__40[23], xbs_fraction__40[24], xbs_fraction__40[25], xbs_fraction__40[26], xbs_fraction__40[27]};
  assign one_hot_159391 = {reverse_159383[27:0] == 28'h000_0000, reverse_159383[27] && reverse_159383[26:0] == 27'h000_0000, reverse_159383[26] && reverse_159383[25:0] == 26'h000_0000, reverse_159383[25] && reverse_159383[24:0] == 25'h000_0000, reverse_159383[24] && reverse_159383[23:0] == 24'h00_0000, reverse_159383[23] && reverse_159383[22:0] == 23'h00_0000, reverse_159383[22] && reverse_159383[21:0] == 22'h00_0000, reverse_159383[21] && reverse_159383[20:0] == 21'h00_0000, reverse_159383[20] && reverse_159383[19:0] == 20'h0_0000, reverse_159383[19] && reverse_159383[18:0] == 19'h0_0000, reverse_159383[18] && reverse_159383[17:0] == 18'h0_0000, reverse_159383[17] && reverse_159383[16:0] == 17'h0_0000, reverse_159383[16] && reverse_159383[15:0] == 16'h0000, reverse_159383[15] && reverse_159383[14:0] == 15'h0000, reverse_159383[14] && reverse_159383[13:0] == 14'h0000, reverse_159383[13] && reverse_159383[12:0] == 13'h0000, reverse_159383[12] && reverse_159383[11:0] == 12'h000, reverse_159383[11] && reverse_159383[10:0] == 11'h000, reverse_159383[10] && reverse_159383[9:0] == 10'h000, reverse_159383[9] && reverse_159383[8:0] == 9'h000, reverse_159383[8] && reverse_159383[7:0] == 8'h00, reverse_159383[7] && reverse_159383[6:0] == 7'h00, reverse_159383[6] && reverse_159383[5:0] == 6'h00, reverse_159383[5] && reverse_159383[4:0] == 5'h00, reverse_159383[4] && reverse_159383[3:0] == 4'h0, reverse_159383[3] && reverse_159383[2:0] == 3'h0, reverse_159383[2] && reverse_159383[1:0] == 2'h0, reverse_159383[1] && !reverse_159383[0], reverse_159383[0]};
  assign reverse_159392 = {xbs_fraction__58[0], xbs_fraction__58[1], xbs_fraction__58[2], xbs_fraction__58[3], xbs_fraction__58[4], xbs_fraction__58[5], xbs_fraction__58[6], xbs_fraction__58[7], xbs_fraction__58[8], xbs_fraction__58[9], xbs_fraction__58[10], xbs_fraction__58[11], xbs_fraction__58[12], xbs_fraction__58[13], xbs_fraction__58[14], xbs_fraction__58[15], xbs_fraction__58[16], xbs_fraction__58[17], xbs_fraction__58[18], xbs_fraction__58[19], xbs_fraction__58[20], xbs_fraction__58[21], xbs_fraction__58[22], xbs_fraction__58[23], xbs_fraction__58[24], xbs_fraction__58[25], xbs_fraction__58[26], xbs_fraction__58[27]};
  assign one_hot_159393 = {reverse_159385[27:0] == 28'h000_0000, reverse_159385[27] && reverse_159385[26:0] == 27'h000_0000, reverse_159385[26] && reverse_159385[25:0] == 26'h000_0000, reverse_159385[25] && reverse_159385[24:0] == 25'h000_0000, reverse_159385[24] && reverse_159385[23:0] == 24'h00_0000, reverse_159385[23] && reverse_159385[22:0] == 23'h00_0000, reverse_159385[22] && reverse_159385[21:0] == 22'h00_0000, reverse_159385[21] && reverse_159385[20:0] == 21'h00_0000, reverse_159385[20] && reverse_159385[19:0] == 20'h0_0000, reverse_159385[19] && reverse_159385[18:0] == 19'h0_0000, reverse_159385[18] && reverse_159385[17:0] == 18'h0_0000, reverse_159385[17] && reverse_159385[16:0] == 17'h0_0000, reverse_159385[16] && reverse_159385[15:0] == 16'h0000, reverse_159385[15] && reverse_159385[14:0] == 15'h0000, reverse_159385[14] && reverse_159385[13:0] == 14'h0000, reverse_159385[13] && reverse_159385[12:0] == 13'h0000, reverse_159385[12] && reverse_159385[11:0] == 12'h000, reverse_159385[11] && reverse_159385[10:0] == 11'h000, reverse_159385[10] && reverse_159385[9:0] == 10'h000, reverse_159385[9] && reverse_159385[8:0] == 9'h000, reverse_159385[8] && reverse_159385[7:0] == 8'h00, reverse_159385[7] && reverse_159385[6:0] == 7'h00, reverse_159385[6] && reverse_159385[5:0] == 6'h00, reverse_159385[5] && reverse_159385[4:0] == 5'h00, reverse_159385[4] && reverse_159385[3:0] == 4'h0, reverse_159385[3] && reverse_159385[2:0] == 3'h0, reverse_159385[2] && reverse_159385[1:0] == 2'h0, reverse_159385[1] && !reverse_159385[0], reverse_159385[0]};
  assign one_hot_159394 = {reverse_159386[27:0] == 28'h000_0000, reverse_159386[27] && reverse_159386[26:0] == 27'h000_0000, reverse_159386[26] && reverse_159386[25:0] == 26'h000_0000, reverse_159386[25] && reverse_159386[24:0] == 25'h000_0000, reverse_159386[24] && reverse_159386[23:0] == 24'h00_0000, reverse_159386[23] && reverse_159386[22:0] == 23'h00_0000, reverse_159386[22] && reverse_159386[21:0] == 22'h00_0000, reverse_159386[21] && reverse_159386[20:0] == 21'h00_0000, reverse_159386[20] && reverse_159386[19:0] == 20'h0_0000, reverse_159386[19] && reverse_159386[18:0] == 19'h0_0000, reverse_159386[18] && reverse_159386[17:0] == 18'h0_0000, reverse_159386[17] && reverse_159386[16:0] == 17'h0_0000, reverse_159386[16] && reverse_159386[15:0] == 16'h0000, reverse_159386[15] && reverse_159386[14:0] == 15'h0000, reverse_159386[14] && reverse_159386[13:0] == 14'h0000, reverse_159386[13] && reverse_159386[12:0] == 13'h0000, reverse_159386[12] && reverse_159386[11:0] == 12'h000, reverse_159386[11] && reverse_159386[10:0] == 11'h000, reverse_159386[10] && reverse_159386[9:0] == 10'h000, reverse_159386[9] && reverse_159386[8:0] == 9'h000, reverse_159386[8] && reverse_159386[7:0] == 8'h00, reverse_159386[7] && reverse_159386[6:0] == 7'h00, reverse_159386[6] && reverse_159386[5:0] == 6'h00, reverse_159386[5] && reverse_159386[4:0] == 5'h00, reverse_159386[4] && reverse_159386[3:0] == 4'h0, reverse_159386[3] && reverse_159386[2:0] == 3'h0, reverse_159386[2] && reverse_159386[1:0] == 2'h0, reverse_159386[1] && !reverse_159386[0], reverse_159386[0]};
  assign encode_159395 = {one_hot_159387[16] | one_hot_159387[17] | one_hot_159387[18] | one_hot_159387[19] | one_hot_159387[20] | one_hot_159387[21] | one_hot_159387[22] | one_hot_159387[23] | one_hot_159387[24] | one_hot_159387[25] | one_hot_159387[26] | one_hot_159387[27] | one_hot_159387[28], one_hot_159387[8] | one_hot_159387[9] | one_hot_159387[10] | one_hot_159387[11] | one_hot_159387[12] | one_hot_159387[13] | one_hot_159387[14] | one_hot_159387[15] | one_hot_159387[24] | one_hot_159387[25] | one_hot_159387[26] | one_hot_159387[27] | one_hot_159387[28], one_hot_159387[4] | one_hot_159387[5] | one_hot_159387[6] | one_hot_159387[7] | one_hot_159387[12] | one_hot_159387[13] | one_hot_159387[14] | one_hot_159387[15] | one_hot_159387[20] | one_hot_159387[21] | one_hot_159387[22] | one_hot_159387[23] | one_hot_159387[28], one_hot_159387[2] | one_hot_159387[3] | one_hot_159387[6] | one_hot_159387[7] | one_hot_159387[10] | one_hot_159387[11] | one_hot_159387[14] | one_hot_159387[15] | one_hot_159387[18] | one_hot_159387[19] | one_hot_159387[22] | one_hot_159387[23] | one_hot_159387[26] | one_hot_159387[27], one_hot_159387[1] | one_hot_159387[3] | one_hot_159387[5] | one_hot_159387[7] | one_hot_159387[9] | one_hot_159387[11] | one_hot_159387[13] | one_hot_159387[15] | one_hot_159387[17] | one_hot_159387[19] | one_hot_159387[21] | one_hot_159387[23] | one_hot_159387[25] | one_hot_159387[27]};
  assign one_hot_159396 = {reverse_159388[27:0] == 28'h000_0000, reverse_159388[27] && reverse_159388[26:0] == 27'h000_0000, reverse_159388[26] && reverse_159388[25:0] == 26'h000_0000, reverse_159388[25] && reverse_159388[24:0] == 25'h000_0000, reverse_159388[24] && reverse_159388[23:0] == 24'h00_0000, reverse_159388[23] && reverse_159388[22:0] == 23'h00_0000, reverse_159388[22] && reverse_159388[21:0] == 22'h00_0000, reverse_159388[21] && reverse_159388[20:0] == 21'h00_0000, reverse_159388[20] && reverse_159388[19:0] == 20'h0_0000, reverse_159388[19] && reverse_159388[18:0] == 19'h0_0000, reverse_159388[18] && reverse_159388[17:0] == 18'h0_0000, reverse_159388[17] && reverse_159388[16:0] == 17'h0_0000, reverse_159388[16] && reverse_159388[15:0] == 16'h0000, reverse_159388[15] && reverse_159388[14:0] == 15'h0000, reverse_159388[14] && reverse_159388[13:0] == 14'h0000, reverse_159388[13] && reverse_159388[12:0] == 13'h0000, reverse_159388[12] && reverse_159388[11:0] == 12'h000, reverse_159388[11] && reverse_159388[10:0] == 11'h000, reverse_159388[10] && reverse_159388[9:0] == 10'h000, reverse_159388[9] && reverse_159388[8:0] == 9'h000, reverse_159388[8] && reverse_159388[7:0] == 8'h00, reverse_159388[7] && reverse_159388[6:0] == 7'h00, reverse_159388[6] && reverse_159388[5:0] == 6'h00, reverse_159388[5] && reverse_159388[4:0] == 5'h00, reverse_159388[4] && reverse_159388[3:0] == 4'h0, reverse_159388[3] && reverse_159388[2:0] == 3'h0, reverse_159388[2] && reverse_159388[1:0] == 2'h0, reverse_159388[1] && !reverse_159388[0], reverse_159388[0]};
  assign encode_159397 = {one_hot_159389[16] | one_hot_159389[17] | one_hot_159389[18] | one_hot_159389[19] | one_hot_159389[20] | one_hot_159389[21] | one_hot_159389[22] | one_hot_159389[23] | one_hot_159389[24] | one_hot_159389[25] | one_hot_159389[26] | one_hot_159389[27] | one_hot_159389[28], one_hot_159389[8] | one_hot_159389[9] | one_hot_159389[10] | one_hot_159389[11] | one_hot_159389[12] | one_hot_159389[13] | one_hot_159389[14] | one_hot_159389[15] | one_hot_159389[24] | one_hot_159389[25] | one_hot_159389[26] | one_hot_159389[27] | one_hot_159389[28], one_hot_159389[4] | one_hot_159389[5] | one_hot_159389[6] | one_hot_159389[7] | one_hot_159389[12] | one_hot_159389[13] | one_hot_159389[14] | one_hot_159389[15] | one_hot_159389[20] | one_hot_159389[21] | one_hot_159389[22] | one_hot_159389[23] | one_hot_159389[28], one_hot_159389[2] | one_hot_159389[3] | one_hot_159389[6] | one_hot_159389[7] | one_hot_159389[10] | one_hot_159389[11] | one_hot_159389[14] | one_hot_159389[15] | one_hot_159389[18] | one_hot_159389[19] | one_hot_159389[22] | one_hot_159389[23] | one_hot_159389[26] | one_hot_159389[27], one_hot_159389[1] | one_hot_159389[3] | one_hot_159389[5] | one_hot_159389[7] | one_hot_159389[9] | one_hot_159389[11] | one_hot_159389[13] | one_hot_159389[15] | one_hot_159389[17] | one_hot_159389[19] | one_hot_159389[21] | one_hot_159389[23] | one_hot_159389[25] | one_hot_159389[27]};
  assign one_hot_159398 = {reverse_159390[27:0] == 28'h000_0000, reverse_159390[27] && reverse_159390[26:0] == 27'h000_0000, reverse_159390[26] && reverse_159390[25:0] == 26'h000_0000, reverse_159390[25] && reverse_159390[24:0] == 25'h000_0000, reverse_159390[24] && reverse_159390[23:0] == 24'h00_0000, reverse_159390[23] && reverse_159390[22:0] == 23'h00_0000, reverse_159390[22] && reverse_159390[21:0] == 22'h00_0000, reverse_159390[21] && reverse_159390[20:0] == 21'h00_0000, reverse_159390[20] && reverse_159390[19:0] == 20'h0_0000, reverse_159390[19] && reverse_159390[18:0] == 19'h0_0000, reverse_159390[18] && reverse_159390[17:0] == 18'h0_0000, reverse_159390[17] && reverse_159390[16:0] == 17'h0_0000, reverse_159390[16] && reverse_159390[15:0] == 16'h0000, reverse_159390[15] && reverse_159390[14:0] == 15'h0000, reverse_159390[14] && reverse_159390[13:0] == 14'h0000, reverse_159390[13] && reverse_159390[12:0] == 13'h0000, reverse_159390[12] && reverse_159390[11:0] == 12'h000, reverse_159390[11] && reverse_159390[10:0] == 11'h000, reverse_159390[10] && reverse_159390[9:0] == 10'h000, reverse_159390[9] && reverse_159390[8:0] == 9'h000, reverse_159390[8] && reverse_159390[7:0] == 8'h00, reverse_159390[7] && reverse_159390[6:0] == 7'h00, reverse_159390[6] && reverse_159390[5:0] == 6'h00, reverse_159390[5] && reverse_159390[4:0] == 5'h00, reverse_159390[4] && reverse_159390[3:0] == 4'h0, reverse_159390[3] && reverse_159390[2:0] == 3'h0, reverse_159390[2] && reverse_159390[1:0] == 2'h0, reverse_159390[1] && !reverse_159390[0], reverse_159390[0]};
  assign encode_159399 = {one_hot_159391[16] | one_hot_159391[17] | one_hot_159391[18] | one_hot_159391[19] | one_hot_159391[20] | one_hot_159391[21] | one_hot_159391[22] | one_hot_159391[23] | one_hot_159391[24] | one_hot_159391[25] | one_hot_159391[26] | one_hot_159391[27] | one_hot_159391[28], one_hot_159391[8] | one_hot_159391[9] | one_hot_159391[10] | one_hot_159391[11] | one_hot_159391[12] | one_hot_159391[13] | one_hot_159391[14] | one_hot_159391[15] | one_hot_159391[24] | one_hot_159391[25] | one_hot_159391[26] | one_hot_159391[27] | one_hot_159391[28], one_hot_159391[4] | one_hot_159391[5] | one_hot_159391[6] | one_hot_159391[7] | one_hot_159391[12] | one_hot_159391[13] | one_hot_159391[14] | one_hot_159391[15] | one_hot_159391[20] | one_hot_159391[21] | one_hot_159391[22] | one_hot_159391[23] | one_hot_159391[28], one_hot_159391[2] | one_hot_159391[3] | one_hot_159391[6] | one_hot_159391[7] | one_hot_159391[10] | one_hot_159391[11] | one_hot_159391[14] | one_hot_159391[15] | one_hot_159391[18] | one_hot_159391[19] | one_hot_159391[22] | one_hot_159391[23] | one_hot_159391[26] | one_hot_159391[27], one_hot_159391[1] | one_hot_159391[3] | one_hot_159391[5] | one_hot_159391[7] | one_hot_159391[9] | one_hot_159391[11] | one_hot_159391[13] | one_hot_159391[15] | one_hot_159391[17] | one_hot_159391[19] | one_hot_159391[21] | one_hot_159391[23] | one_hot_159391[25] | one_hot_159391[27]};
  assign one_hot_159400 = {reverse_159392[27:0] == 28'h000_0000, reverse_159392[27] && reverse_159392[26:0] == 27'h000_0000, reverse_159392[26] && reverse_159392[25:0] == 26'h000_0000, reverse_159392[25] && reverse_159392[24:0] == 25'h000_0000, reverse_159392[24] && reverse_159392[23:0] == 24'h00_0000, reverse_159392[23] && reverse_159392[22:0] == 23'h00_0000, reverse_159392[22] && reverse_159392[21:0] == 22'h00_0000, reverse_159392[21] && reverse_159392[20:0] == 21'h00_0000, reverse_159392[20] && reverse_159392[19:0] == 20'h0_0000, reverse_159392[19] && reverse_159392[18:0] == 19'h0_0000, reverse_159392[18] && reverse_159392[17:0] == 18'h0_0000, reverse_159392[17] && reverse_159392[16:0] == 17'h0_0000, reverse_159392[16] && reverse_159392[15:0] == 16'h0000, reverse_159392[15] && reverse_159392[14:0] == 15'h0000, reverse_159392[14] && reverse_159392[13:0] == 14'h0000, reverse_159392[13] && reverse_159392[12:0] == 13'h0000, reverse_159392[12] && reverse_159392[11:0] == 12'h000, reverse_159392[11] && reverse_159392[10:0] == 11'h000, reverse_159392[10] && reverse_159392[9:0] == 10'h000, reverse_159392[9] && reverse_159392[8:0] == 9'h000, reverse_159392[8] && reverse_159392[7:0] == 8'h00, reverse_159392[7] && reverse_159392[6:0] == 7'h00, reverse_159392[6] && reverse_159392[5:0] == 6'h00, reverse_159392[5] && reverse_159392[4:0] == 5'h00, reverse_159392[4] && reverse_159392[3:0] == 4'h0, reverse_159392[3] && reverse_159392[2:0] == 3'h0, reverse_159392[2] && reverse_159392[1:0] == 2'h0, reverse_159392[1] && !reverse_159392[0], reverse_159392[0]};
  assign encode_159401 = {one_hot_159393[16] | one_hot_159393[17] | one_hot_159393[18] | one_hot_159393[19] | one_hot_159393[20] | one_hot_159393[21] | one_hot_159393[22] | one_hot_159393[23] | one_hot_159393[24] | one_hot_159393[25] | one_hot_159393[26] | one_hot_159393[27] | one_hot_159393[28], one_hot_159393[8] | one_hot_159393[9] | one_hot_159393[10] | one_hot_159393[11] | one_hot_159393[12] | one_hot_159393[13] | one_hot_159393[14] | one_hot_159393[15] | one_hot_159393[24] | one_hot_159393[25] | one_hot_159393[26] | one_hot_159393[27] | one_hot_159393[28], one_hot_159393[4] | one_hot_159393[5] | one_hot_159393[6] | one_hot_159393[7] | one_hot_159393[12] | one_hot_159393[13] | one_hot_159393[14] | one_hot_159393[15] | one_hot_159393[20] | one_hot_159393[21] | one_hot_159393[22] | one_hot_159393[23] | one_hot_159393[28], one_hot_159393[2] | one_hot_159393[3] | one_hot_159393[6] | one_hot_159393[7] | one_hot_159393[10] | one_hot_159393[11] | one_hot_159393[14] | one_hot_159393[15] | one_hot_159393[18] | one_hot_159393[19] | one_hot_159393[22] | one_hot_159393[23] | one_hot_159393[26] | one_hot_159393[27], one_hot_159393[1] | one_hot_159393[3] | one_hot_159393[5] | one_hot_159393[7] | one_hot_159393[9] | one_hot_159393[11] | one_hot_159393[13] | one_hot_159393[15] | one_hot_159393[17] | one_hot_159393[19] | one_hot_159393[21] | one_hot_159393[23] | one_hot_159393[25] | one_hot_159393[27]};
  assign encode_159402 = {one_hot_159394[16] | one_hot_159394[17] | one_hot_159394[18] | one_hot_159394[19] | one_hot_159394[20] | one_hot_159394[21] | one_hot_159394[22] | one_hot_159394[23] | one_hot_159394[24] | one_hot_159394[25] | one_hot_159394[26] | one_hot_159394[27] | one_hot_159394[28], one_hot_159394[8] | one_hot_159394[9] | one_hot_159394[10] | one_hot_159394[11] | one_hot_159394[12] | one_hot_159394[13] | one_hot_159394[14] | one_hot_159394[15] | one_hot_159394[24] | one_hot_159394[25] | one_hot_159394[26] | one_hot_159394[27] | one_hot_159394[28], one_hot_159394[4] | one_hot_159394[5] | one_hot_159394[6] | one_hot_159394[7] | one_hot_159394[12] | one_hot_159394[13] | one_hot_159394[14] | one_hot_159394[15] | one_hot_159394[20] | one_hot_159394[21] | one_hot_159394[22] | one_hot_159394[23] | one_hot_159394[28], one_hot_159394[2] | one_hot_159394[3] | one_hot_159394[6] | one_hot_159394[7] | one_hot_159394[10] | one_hot_159394[11] | one_hot_159394[14] | one_hot_159394[15] | one_hot_159394[18] | one_hot_159394[19] | one_hot_159394[22] | one_hot_159394[23] | one_hot_159394[26] | one_hot_159394[27], one_hot_159394[1] | one_hot_159394[3] | one_hot_159394[5] | one_hot_159394[7] | one_hot_159394[9] | one_hot_159394[11] | one_hot_159394[13] | one_hot_159394[15] | one_hot_159394[17] | one_hot_159394[19] | one_hot_159394[21] | one_hot_159394[23] | one_hot_159394[25] | one_hot_159394[27]};
  assign encode_159404 = {one_hot_159396[16] | one_hot_159396[17] | one_hot_159396[18] | one_hot_159396[19] | one_hot_159396[20] | one_hot_159396[21] | one_hot_159396[22] | one_hot_159396[23] | one_hot_159396[24] | one_hot_159396[25] | one_hot_159396[26] | one_hot_159396[27] | one_hot_159396[28], one_hot_159396[8] | one_hot_159396[9] | one_hot_159396[10] | one_hot_159396[11] | one_hot_159396[12] | one_hot_159396[13] | one_hot_159396[14] | one_hot_159396[15] | one_hot_159396[24] | one_hot_159396[25] | one_hot_159396[26] | one_hot_159396[27] | one_hot_159396[28], one_hot_159396[4] | one_hot_159396[5] | one_hot_159396[6] | one_hot_159396[7] | one_hot_159396[12] | one_hot_159396[13] | one_hot_159396[14] | one_hot_159396[15] | one_hot_159396[20] | one_hot_159396[21] | one_hot_159396[22] | one_hot_159396[23] | one_hot_159396[28], one_hot_159396[2] | one_hot_159396[3] | one_hot_159396[6] | one_hot_159396[7] | one_hot_159396[10] | one_hot_159396[11] | one_hot_159396[14] | one_hot_159396[15] | one_hot_159396[18] | one_hot_159396[19] | one_hot_159396[22] | one_hot_159396[23] | one_hot_159396[26] | one_hot_159396[27], one_hot_159396[1] | one_hot_159396[3] | one_hot_159396[5] | one_hot_159396[7] | one_hot_159396[9] | one_hot_159396[11] | one_hot_159396[13] | one_hot_159396[15] | one_hot_159396[17] | one_hot_159396[19] | one_hot_159396[21] | one_hot_159396[23] | one_hot_159396[25] | one_hot_159396[27]};
  assign encode_159406 = {one_hot_159398[16] | one_hot_159398[17] | one_hot_159398[18] | one_hot_159398[19] | one_hot_159398[20] | one_hot_159398[21] | one_hot_159398[22] | one_hot_159398[23] | one_hot_159398[24] | one_hot_159398[25] | one_hot_159398[26] | one_hot_159398[27] | one_hot_159398[28], one_hot_159398[8] | one_hot_159398[9] | one_hot_159398[10] | one_hot_159398[11] | one_hot_159398[12] | one_hot_159398[13] | one_hot_159398[14] | one_hot_159398[15] | one_hot_159398[24] | one_hot_159398[25] | one_hot_159398[26] | one_hot_159398[27] | one_hot_159398[28], one_hot_159398[4] | one_hot_159398[5] | one_hot_159398[6] | one_hot_159398[7] | one_hot_159398[12] | one_hot_159398[13] | one_hot_159398[14] | one_hot_159398[15] | one_hot_159398[20] | one_hot_159398[21] | one_hot_159398[22] | one_hot_159398[23] | one_hot_159398[28], one_hot_159398[2] | one_hot_159398[3] | one_hot_159398[6] | one_hot_159398[7] | one_hot_159398[10] | one_hot_159398[11] | one_hot_159398[14] | one_hot_159398[15] | one_hot_159398[18] | one_hot_159398[19] | one_hot_159398[22] | one_hot_159398[23] | one_hot_159398[26] | one_hot_159398[27], one_hot_159398[1] | one_hot_159398[3] | one_hot_159398[5] | one_hot_159398[7] | one_hot_159398[9] | one_hot_159398[11] | one_hot_159398[13] | one_hot_159398[15] | one_hot_159398[17] | one_hot_159398[19] | one_hot_159398[21] | one_hot_159398[23] | one_hot_159398[25] | one_hot_159398[27]};
  assign encode_159408 = {one_hot_159400[16] | one_hot_159400[17] | one_hot_159400[18] | one_hot_159400[19] | one_hot_159400[20] | one_hot_159400[21] | one_hot_159400[22] | one_hot_159400[23] | one_hot_159400[24] | one_hot_159400[25] | one_hot_159400[26] | one_hot_159400[27] | one_hot_159400[28], one_hot_159400[8] | one_hot_159400[9] | one_hot_159400[10] | one_hot_159400[11] | one_hot_159400[12] | one_hot_159400[13] | one_hot_159400[14] | one_hot_159400[15] | one_hot_159400[24] | one_hot_159400[25] | one_hot_159400[26] | one_hot_159400[27] | one_hot_159400[28], one_hot_159400[4] | one_hot_159400[5] | one_hot_159400[6] | one_hot_159400[7] | one_hot_159400[12] | one_hot_159400[13] | one_hot_159400[14] | one_hot_159400[15] | one_hot_159400[20] | one_hot_159400[21] | one_hot_159400[22] | one_hot_159400[23] | one_hot_159400[28], one_hot_159400[2] | one_hot_159400[3] | one_hot_159400[6] | one_hot_159400[7] | one_hot_159400[10] | one_hot_159400[11] | one_hot_159400[14] | one_hot_159400[15] | one_hot_159400[18] | one_hot_159400[19] | one_hot_159400[22] | one_hot_159400[23] | one_hot_159400[26] | one_hot_159400[27], one_hot_159400[1] | one_hot_159400[3] | one_hot_159400[5] | one_hot_159400[7] | one_hot_159400[9] | one_hot_159400[11] | one_hot_159400[13] | one_hot_159400[15] | one_hot_159400[17] | one_hot_159400[19] | one_hot_159400[21] | one_hot_159400[23] | one_hot_159400[25] | one_hot_159400[27]};
  assign cancel__11 = |encode_159395[4:1];
  assign carry_bit__10 = xbs_fraction__10[27];
  assign result_fraction__484 = 23'h00_0000;
  assign cancel__22 = |encode_159397[4:1];
  assign carry_bit__22 = xbs_fraction__21[27];
  assign result_fraction__549 = 23'h00_0000;
  assign cancel__41 = |encode_159399[4:1];
  assign carry_bit__41 = xbs_fraction__39[27];
  assign result_fraction__614 = 23'h00_0000;
  assign cancel__60 = |encode_159401[4:1];
  assign carry_bit__60 = xbs_fraction__57[27];
  assign result_fraction__683 = 23'h00_0000;
  assign cancel__1 = |encode_159402[4:1];
  assign carry_bit__2 = xbs_fraction__2[27];
  assign result_fraction__485 = 23'h00_0000;
  assign leading_zeroes__10 = {result_fraction__484, encode_159395};
  assign cancel__23 = |encode_159404[4:1];
  assign carry_bit__23 = xbs_fraction__22[27];
  assign result_fraction__550 = 23'h00_0000;
  assign leading_zeroes__22 = {result_fraction__549, encode_159397};
  assign cancel__42 = |encode_159406[4:1];
  assign carry_bit__42 = xbs_fraction__40[27];
  assign result_fraction__615 = 23'h00_0000;
  assign leading_zeroes__41 = {result_fraction__614, encode_159399};
  assign cancel__61 = |encode_159408[4:1];
  assign carry_bit__61 = xbs_fraction__58[27];
  assign result_fraction__684 = 23'h00_0000;
  assign leading_zeroes__60 = {result_fraction__683, encode_159401};
  assign leading_zeroes__2 = {result_fraction__485, encode_159402};
  assign carry_fraction__20 = xbs_fraction__10[27:1];
  assign add_159476 = leading_zeroes__10 + 28'hfff_ffff;
  assign leading_zeroes__23 = {result_fraction__550, encode_159404};
  assign carry_fraction__43 = xbs_fraction__21[27:1];
  assign add_159489 = leading_zeroes__22 + 28'hfff_ffff;
  assign array_index_159490 = in_img_unflattened[4'h3];
  assign leading_zeroes__42 = {result_fraction__615, encode_159406};
  assign carry_fraction__81 = xbs_fraction__39[27:1];
  assign add_159503 = leading_zeroes__41 + 28'hfff_ffff;
  assign leading_zeroes__61 = {result_fraction__684, encode_159408};
  assign carry_fraction__119 = xbs_fraction__57[27:1];
  assign add_159516 = leading_zeroes__60 + 28'hfff_ffff;
  assign array_index_159517 = in_img_unflattened[4'h7];
  assign carry_fraction__3 = xbs_fraction__2[27:1];
  assign add_159524 = leading_zeroes__2 + 28'hfff_ffff;
  assign concat_159525 = {~(carry_bit__10 | cancel__11), ~(carry_bit__10 | ~cancel__11), ~(~carry_bit__10 | cancel__11)};
  assign carry_fraction__21 = carry_fraction__20 | {26'h000_0000, xbs_fraction__10[0]};
  assign cancel_fraction__10 = add_159476 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__10[26:0] << add_159476;
  assign result_sign__485 = 1'h0;
  assign carry_fraction__44 = xbs_fraction__22[27:1];
  assign add_159535 = leading_zeroes__23 + 28'hfff_ffff;
  assign concat_159536 = {~(carry_bit__22 | cancel__22), ~(carry_bit__22 | ~cancel__22), ~(~carry_bit__22 | cancel__22)};
  assign carry_fraction__45 = carry_fraction__43 | {26'h000_0000, xbs_fraction__21[0]};
  assign cancel_fraction__22 = add_159489 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__21[26:0] << add_159489;
  assign result_sign__492 = 1'h0;
  assign x_bexp__173 = array_index_159490[30:23];
  assign carry_fraction__82 = xbs_fraction__40[27:1];
  assign add_159547 = leading_zeroes__42 + 28'hfff_ffff;
  assign concat_159548 = {~(carry_bit__41 | cancel__41), ~(carry_bit__41 | ~cancel__41), ~(~carry_bit__41 | cancel__41)};
  assign carry_fraction__83 = carry_fraction__81 | {26'h000_0000, xbs_fraction__39[0]};
  assign cancel_fraction__41 = add_159503 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__39[26:0] << add_159503;
  assign result_sign__684 = 1'h0;
  assign carry_fraction__120 = xbs_fraction__58[27:1];
  assign add_159558 = leading_zeroes__61 + 28'hfff_ffff;
  assign concat_159559 = {~(carry_bit__60 | cancel__60), ~(carry_bit__60 | ~cancel__60), ~(~carry_bit__60 | cancel__60)};
  assign carry_fraction__121 = carry_fraction__119 | {26'h000_0000, xbs_fraction__57[0]};
  assign cancel_fraction__60 = add_159516 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__57[26:0] << add_159516;
  assign result_sign__691 = 1'h0;
  assign x_bexp__461 = array_index_159517[30:23];
  assign concat_159564 = {~(carry_bit__2 | cancel__1), ~(carry_bit__2 | ~cancel__1), ~(~carry_bit__2 | cancel__1)};
  assign carry_fraction__4 = carry_fraction__3 | {26'h000_0000, xbs_fraction__2[0]};
  assign cancel_fraction__2 = add_159524 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__2[26:0] << add_159524;
  assign shifted_fraction__10 = carry_fraction__21 & {27{concat_159525[0]}} | cancel_fraction__10 & {27{concat_159525[1]}} | xbs_fraction__10[26:0] & {27{concat_159525[2]}};
  assign concat_159570 = {~(carry_bit__23 | cancel__23), ~(carry_bit__23 | ~cancel__23), ~(~carry_bit__23 | cancel__23)};
  assign carry_fraction__46 = carry_fraction__44 | {26'h000_0000, xbs_fraction__22[0]};
  assign cancel_fraction__23 = add_159535 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__22[26:0] << add_159535;
  assign shifted_fraction__22 = carry_fraction__45 & {27{concat_159536[0]}} | cancel_fraction__22 & {27{concat_159536[1]}} | xbs_fraction__21[26:0] & {27{concat_159536[2]}};
  assign concat_159576 = {~(carry_bit__42 | cancel__42), ~(carry_bit__42 | ~cancel__42), ~(~carry_bit__42 | cancel__42)};
  assign carry_fraction__84 = carry_fraction__82 | {26'h000_0000, xbs_fraction__40[0]};
  assign cancel_fraction__42 = add_159547 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__40[26:0] << add_159547;
  assign shifted_fraction__41 = carry_fraction__83 & {27{concat_159548[0]}} | cancel_fraction__41 & {27{concat_159548[1]}} | xbs_fraction__39[26:0] & {27{concat_159548[2]}};
  assign concat_159582 = {~(carry_bit__61 | cancel__61), ~(carry_bit__61 | ~cancel__61), ~(~carry_bit__61 | cancel__61)};
  assign carry_fraction__122 = carry_fraction__120 | {26'h000_0000, xbs_fraction__58[0]};
  assign cancel_fraction__61 = add_159558 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__58[26:0] << add_159558;
  assign shifted_fraction__60 = carry_fraction__121 & {27{concat_159559[0]}} | cancel_fraction__60 & {27{concat_159559[1]}} | xbs_fraction__57[26:0] & {27{concat_159559[2]}};
  assign shifted_fraction__2 = carry_fraction__4 & {27{concat_159564[0]}} | cancel_fraction__2 & {27{concat_159564[1]}} | xbs_fraction__2[26:0] & {27{concat_159564[2]}};
  assign result_sign__972 = 1'h0;
  assign result_sign__398 = 1'h0;
  assign add_159592 = {result_sign__485, x_bexp__157} + 9'h07f;
  assign shifted_fraction__23 = carry_fraction__46 & {27{concat_159570[0]}} | cancel_fraction__23 & {27{concat_159570[1]}} | xbs_fraction__22[26:0] & {27{concat_159570[2]}};
  assign result_sign__973 = 1'h0;
  assign result_sign__495 = 1'h0;
  assign add_159597 = {result_sign__492, x_bexp__173} + 9'h07f;
  assign x_bexp__690 = 8'h00;
  assign result_sign__491 = 1'h0;
  assign x_fraction__173 = array_index_159490[22:0];
  assign shifted_fraction__42 = carry_fraction__84 & {27{concat_159576[0]}} | cancel_fraction__42 & {27{concat_159576[1]}} | xbs_fraction__40[26:0] & {27{concat_159576[2]}};
  assign result_sign__974 = 1'h0;
  assign result_sign__588 = 1'h0;
  assign add_159605 = {result_sign__684, x_bexp__445} + 9'h07f;
  assign shifted_fraction__61 = carry_fraction__122 & {27{concat_159582[0]}} | cancel_fraction__61 & {27{concat_159582[1]}} | xbs_fraction__58[26:0] & {27{concat_159582[2]}};
  assign result_sign__975 = 1'h0;
  assign result_sign__694 = 1'h0;
  assign add_159610 = {result_sign__691, x_bexp__461} + 9'h07f;
  assign x_bexp__691 = 8'h00;
  assign result_sign__690 = 1'h0;
  assign x_fraction__461 = array_index_159517[22:0];
  assign result_sign__976 = 1'h0;
  assign normal_chunk__10 = shifted_fraction__10[2:0];
  assign fraction_shift__229 = 3'h4;
  assign half_way_chunk__10 = shifted_fraction__10[3:2];
  assign result_sign__977 = 1'h0;
  assign normal_chunk__22 = shifted_fraction__22[2:0];
  assign fraction_shift__264 = 3'h4;
  assign half_way_chunk__22 = shifted_fraction__22[3:2];
  assign ne_159634 = x_bexp__173 != x_bexp__690;
  assign result_sign__978 = 1'h0;
  assign normal_chunk__41 = shifted_fraction__41[2:0];
  assign fraction_shift__299 = 3'h4;
  assign half_way_chunk__41 = shifted_fraction__41[3:2];
  assign result_sign__979 = 1'h0;
  assign normal_chunk__60 = shifted_fraction__60[2:0];
  assign fraction_shift__334 = 3'h4;
  assign half_way_chunk__60 = shifted_fraction__60[3:2];
  assign ne_159657 = x_bexp__461 != x_bexp__691;
  assign normal_chunk__2 = shifted_fraction__2[2:0];
  assign fraction_shift__230 = 3'h4;
  assign half_way_chunk__2 = shifted_fraction__2[3:2];
  assign result_sign__396 = 1'h0;
  assign add_159669 = {result_sign__972, shifted_fraction__10[26:3]} + 25'h000_0001;
  assign exp__44 = {result_sign__398, add_159592} + 10'h381;
  assign normal_chunk__23 = shifted_fraction__23[2:0];
  assign fraction_shift__265 = 3'h4;
  assign half_way_chunk__23 = shifted_fraction__23[3:2];
  assign result_sign__493 = 1'h0;
  assign add_159680 = {result_sign__973, shifted_fraction__22[26:3]} + 25'h000_0001;
  assign exp__99 = {result_sign__495, add_159597} + 10'h381;
  assign x_fraction__175 = {result_sign__491, x_fraction__173} | 24'h80_0000;
  assign normal_chunk__42 = shifted_fraction__42[2:0];
  assign fraction_shift__300 = 3'h4;
  assign half_way_chunk__42 = shifted_fraction__42[3:2];
  assign result_sign__586 = 1'h0;
  assign add_159694 = {result_sign__974, shifted_fraction__41[26:3]} + 25'h000_0001;
  assign exp__181 = {result_sign__588, add_159605} + 10'h381;
  assign normal_chunk__61 = shifted_fraction__61[2:0];
  assign fraction_shift__335 = 3'h4;
  assign half_way_chunk__61 = shifted_fraction__61[3:2];
  assign result_sign__692 = 1'h0;
  assign add_159705 = {result_sign__975, shifted_fraction__60[26:3]} + 25'h000_0001;
  assign exp__263 = {result_sign__694, add_159610} + 10'h381;
  assign sign_ext_159707 = {10{ne_159657}};
  assign x_fraction__463 = {result_sign__690, x_fraction__461} | 24'h80_0000;
  assign result_sign__397 = 1'h0;
  assign add_159713 = {result_sign__976, shifted_fraction__2[26:3]} + 25'h000_0001;
  assign do_round_up__21 = normal_chunk__10 > fraction_shift__229 | half_way_chunk__10 == 2'h3;
  assign exp__45 = exp__44 & sign_ext_158460;
  assign result_sign__494 = 1'h0;
  assign add_159722 = {result_sign__977, shifted_fraction__23[26:3]} + 25'h000_0001;
  assign do_round_up__46 = normal_chunk__22 > fraction_shift__264 | half_way_chunk__22 == 2'h3;
  assign exp__101 = exp__99 & {10{ne_159634}};
  assign x_fraction__177 = x_fraction__175 & {24{ne_159634}};
  assign result_sign__808 = 1'h0;
  assign result_sign__809 = 1'h0;
  assign result_sign__587 = 1'h0;
  assign add_159734 = {result_sign__978, shifted_fraction__42[26:3]} + 25'h000_0001;
  assign do_round_up__85 = normal_chunk__41 > fraction_shift__299 | half_way_chunk__41 == 2'h3;
  assign exp__183 = exp__181 & sign_ext_158473;
  assign result_sign__693 = 1'h0;
  assign add_159743 = {result_sign__979, shifted_fraction__61[26:3]} + 25'h000_0001;
  assign do_round_up__124 = normal_chunk__60 > fraction_shift__334 | half_way_chunk__60 == 2'h3;
  assign exp__265 = exp__263 & sign_ext_159707;
  assign x_fraction__465 = x_fraction__463 & {24{ne_159657}};
  assign result_sign__810 = 1'h0;
  assign result_sign__811 = 1'h0;
  assign do_round_up__4 = normal_chunk__2 > fraction_shift__230 | half_way_chunk__2 == 2'h3;
  assign rounded_fraction__10 = do_round_up__21 ? {add_159669, normal_chunk__10} : {result_sign__396, shifted_fraction__10};
  assign do_round_up__47 = normal_chunk__23 > fraction_shift__265 | half_way_chunk__23 == 2'h3;
  assign rounded_fraction__22 = do_round_up__46 ? {add_159680, normal_chunk__22} : {result_sign__493, shifted_fraction__22};
  assign do_round_up__86 = normal_chunk__42 > fraction_shift__300 | half_way_chunk__42 == 2'h3;
  assign rounded_fraction__41 = do_round_up__85 ? {add_159694, normal_chunk__41} : {result_sign__586, shifted_fraction__41};
  assign do_round_up__125 = normal_chunk__61 > fraction_shift__335 | half_way_chunk__61 == 2'h3;
  assign rounded_fraction__60 = do_round_up__124 ? {add_159705, normal_chunk__60} : {result_sign__692, shifted_fraction__60};
  assign concat_159774 = {x_fraction__465, result_sign__810};
  assign concat_159775 = {result_sign__811, x_fraction__465};
  assign rounded_fraction__2 = do_round_up__4 ? {add_159713, normal_chunk__2} : {result_sign__397, shifted_fraction__2};
  assign result_sign__399 = 1'h0;
  assign x_bexp__77 = 8'h00;
  assign rounding_carry__10 = rounded_fraction__10[27];
  assign sel_159780 = $signed(exp__45) <= $signed(10'h000) ? concat_158507 : concat_158506;
  assign rounded_fraction__23 = do_round_up__47 ? {add_159722, normal_chunk__23} : {result_sign__494, shifted_fraction__23};
  assign result_sign__496 = 1'h0;
  assign x_bexp__594 = 8'h00;
  assign rounding_carry__22 = rounded_fraction__22[27];
  assign sel_159785 = $signed(exp__101) <= $signed(10'h000) ? {result_sign__809, x_fraction__177} : {x_fraction__177, result_sign__808};
  assign rounded_fraction__42 = do_round_up__86 ? {add_159734, normal_chunk__42} : {result_sign__587, shifted_fraction__42};
  assign result_sign__589 = 1'h0;
  assign x_bexp__612 = 8'h00;
  assign rounding_carry__41 = rounded_fraction__41[27];
  assign sel_159790 = $signed(exp__183) <= $signed(10'h000) ? concat_158513 : concat_158512;
  assign rounded_fraction__61 = do_round_up__125 ? {add_159743, normal_chunk__61} : {result_sign__693, shifted_fraction__61};
  assign result_sign__695 = 1'h0;
  assign x_bexp__630 = 8'h00;
  assign rounding_carry__60 = rounded_fraction__60[27];
  assign sel_159795 = $signed(exp__265) <= $signed(10'h000) ? concat_159775 : concat_159774;
  assign result_sign__400 = 1'h0;
  assign x_bexp__577 = 8'h00;
  assign rounding_carry__2 = rounded_fraction__2[27];
  assign result_sign__930 = 1'h0;
  assign fraction__104 = sel_159780[23:1];
  assign result_sign__497 = 1'h0;
  assign x_bexp__595 = 8'h00;
  assign rounding_carry__23 = rounded_fraction__23[27];
  assign result_sign__936 = 1'h0;
  assign fraction__226 = sel_159785[23:1];
  assign result_sign__590 = 1'h0;
  assign x_bexp__613 = 8'h00;
  assign rounding_carry__42 = rounded_fraction__42[27];
  assign result_sign__942 = 1'h0;
  assign fraction__405 = sel_159790[23:1];
  assign result_sign__696 = 1'h0;
  assign x_bexp__631 = 8'h00;
  assign rounding_carry__61 = rounded_fraction__61[27];
  assign result_sign__950 = 1'h0;
  assign fraction__584 = sel_159795[23:1];
  assign result_sign__401 = 1'h0;
  assign add_159827 = {result_sign__399, x_bexp__86} + {x_bexp__77, rounding_carry__10};
  assign fraction__105 = {result_sign__930, fraction__104};
  assign result_sign__498 = 1'h0;
  assign add_159837 = {result_sign__496, x_bexp__171} + {x_bexp__594, rounding_carry__22};
  assign fraction__228 = {result_sign__936, fraction__226};
  assign result_sign__591 = 1'h0;
  assign add_159847 = {result_sign__589, x_bexp__315} + {x_bexp__612, rounding_carry__41};
  assign fraction__407 = {result_sign__942, fraction__405};
  assign result_sign__697 = 1'h0;
  assign add_159857 = {result_sign__695, x_bexp__459} + {x_bexp__630, rounding_carry__60};
  assign fraction__586 = {result_sign__950, fraction__584};
  assign result_sign__402 = 1'h0;
  assign add_159865 = {result_sign__400, x_bexp__14} + {x_bexp__577, rounding_carry__2};
  assign do_round_up__22 = sel_159780[0] & sel_159780[1];
  assign add_159874 = fraction__105 + 24'h00_0001;
  assign result_sign__499 = 1'h0;
  assign add_159876 = {result_sign__497, x_bexp__172} + {x_bexp__595, rounding_carry__23};
  assign do_round_up__48 = sel_159785[0] & sel_159785[1];
  assign add_159885 = fraction__228 + 24'h00_0001;
  assign result_sign__592 = 1'h0;
  assign add_159887 = {result_sign__590, x_bexp__316} + {x_bexp__613, rounding_carry__42};
  assign do_round_up__87 = sel_159790[0] & sel_159790[1];
  assign add_159896 = fraction__407 + 24'h00_0001;
  assign result_sign__698 = 1'h0;
  assign add_159898 = {result_sign__696, x_bexp__460} + {x_bexp__631, rounding_carry__61};
  assign do_round_up__126 = sel_159795[0] & sel_159795[1];
  assign add_159907 = fraction__586 + 24'h00_0001;
  assign add_159913 = {result_sign__401, add_159827} + 10'h001;
  assign fraction__106 = do_round_up__22 ? add_159874 : fraction__105;
  assign add_159923 = {result_sign__498, add_159837} + 10'h001;
  assign fraction__230 = do_round_up__48 ? add_159885 : fraction__228;
  assign add_159933 = {result_sign__591, add_159847} + 10'h001;
  assign fraction__409 = do_round_up__87 ? add_159896 : fraction__407;
  assign add_159943 = {result_sign__697, add_159857} + 10'h001;
  assign fraction__588 = do_round_up__126 ? add_159907 : fraction__586;
  assign add_159948 = {result_sign__402, add_159865} + 10'h001;
  assign wide_exponent__30 = add_159913 - {5'h00, encode_159395};
  assign add_159954 = exp__45 + 10'h001;
  assign add_159955 = {result_sign__499, add_159876} + 10'h001;
  assign wide_exponent__64 = add_159923 - {5'h00, encode_159397};
  assign add_159961 = exp__101 + 10'h001;
  assign add_159962 = {result_sign__592, add_159887} + 10'h001;
  assign wide_exponent__121 = add_159933 - {5'h00, encode_159399};
  assign add_159968 = exp__183 + 10'h001;
  assign add_159969 = {result_sign__698, add_159898} + 10'h001;
  assign wide_exponent__178 = add_159943 - {5'h00, encode_159401};
  assign add_159975 = exp__265 + 10'h001;
  assign wide_exponent__4 = add_159948 - {5'h00, encode_159402};
  assign wide_exponent__31 = wide_exponent__30 & {10{add_159320 != 26'h000_0000 | xddend_y__10[2:0] != 3'h0}};
  assign exp__47 = fraction__106[23] ? add_159954 : exp__45;
  assign wide_exponent__65 = add_159955 - {5'h00, encode_159404};
  assign wide_exponent__66 = wide_exponent__64 & {10{add_159323 != 26'h000_0000 | xddend_y__21[2:0] != 3'h0}};
  assign exp__105 = fraction__230[23] ? add_159961 : exp__101;
  assign wide_exponent__122 = add_159962 - {5'h00, encode_159406};
  assign wide_exponent__123 = wide_exponent__121 & {10{add_159326 != 26'h000_0000 | xddend_y__39[2:0] != 3'h0}};
  assign exp__187 = fraction__409[23] ? add_159968 : exp__183;
  assign wide_exponent__179 = add_159969 - {5'h00, encode_159408};
  assign wide_exponent__180 = wide_exponent__178 & {10{add_159329 != 26'h000_0000 | xddend_y__57[2:0] != 3'h0}};
  assign exp__269 = fraction__588[23] ? add_159975 : exp__265;
  assign wide_exponent__5 = wide_exponent__4 & {10{add_159330 != 26'h000_0000 | xddend_y__2[2:0] != 3'h0}};
  assign high_exp__365 = 8'hff;
  assign result_fraction__771 = 23'h00_0000;
  assign high_exp__366 = 8'hff;
  assign result_fraction__772 = 23'h00_0000;
  assign high_exp__84 = 8'hff;
  assign result_fraction__486 = 23'h00_0000;
  assign high_exp__85 = 8'hff;
  assign result_fraction__487 = 23'h00_0000;
  assign wide_exponent__67 = wide_exponent__65 & {10{add_159333 != 26'h000_0000 | xddend_y__22[2:0] != 3'h0}};
  assign high_exp__397 = 8'hff;
  assign result_fraction__804 = 23'h00_0000;
  assign high_exp__398 = 8'hff;
  assign result_fraction__805 = 23'h00_0000;
  assign high_exp__148 = 8'hff;
  assign result_fraction__551 = 23'h00_0000;
  assign high_exp__149 = 8'hff;
  assign result_fraction__552 = 23'h00_0000;
  assign wide_exponent__124 = wide_exponent__122 & {10{add_159336 != 26'h000_0000 | xddend_y__40[2:0] != 3'h0}};
  assign high_exp__429 = 8'hff;
  assign result_fraction__837 = 23'h00_0000;
  assign high_exp__430 = 8'hff;
  assign result_fraction__838 = 23'h00_0000;
  assign high_exp__213 = 8'hff;
  assign result_fraction__616 = 23'h00_0000;
  assign high_exp__214 = 8'hff;
  assign result_fraction__617 = 23'h00_0000;
  assign wide_exponent__181 = wide_exponent__179 & {10{add_159339 != 26'h000_0000 | xddend_y__58[2:0] != 3'h0}};
  assign high_exp__461 = 8'hff;
  assign result_fraction__870 = 23'h00_0000;
  assign high_exp__462 = 8'hff;
  assign result_fraction__871 = 23'h00_0000;
  assign high_exp__282 = 8'hff;
  assign result_fraction__685 = 23'h00_0000;
  assign high_exp__283 = 8'hff;
  assign result_fraction__686 = 23'h00_0000;
  assign ne_160043 = x_fraction__86 != result_fraction__771;
  assign ne_160045 = prod_fraction__30 != result_fraction__772;
  assign eq_160046 = x_bexp__86 == high_exp__84;
  assign eq_160047 = x_fraction__86 == result_fraction__486;
  assign eq_160048 = prod_bexp__42 == high_exp__85;
  assign eq_160049 = prod_fraction__30 == result_fraction__487;
  assign result_exp__33 = exp__47[8:0];
  assign ne_160055 = x_fraction__171 != result_fraction__804;
  assign ne_160057 = prod_fraction__61 != result_fraction__805;
  assign eq_160058 = x_bexp__171 == high_exp__148;
  assign eq_160059 = x_fraction__171 == result_fraction__551;
  assign eq_160060 = prod_bexp__83 == high_exp__149;
  assign eq_160061 = prod_fraction__61 == result_fraction__552;
  assign result_exp__73 = exp__105[8:0];
  assign ne_160067 = x_fraction__315 != result_fraction__837;
  assign ne_160069 = prod_fraction__115 != result_fraction__838;
  assign eq_160070 = x_bexp__315 == high_exp__213;
  assign eq_160071 = x_fraction__315 == result_fraction__616;
  assign eq_160072 = prod_bexp__155 == high_exp__214;
  assign eq_160073 = prod_fraction__115 == result_fraction__617;
  assign result_exp__133 = exp__187[8:0];
  assign ne_160079 = x_fraction__459 != result_fraction__870;
  assign ne_160081 = prod_fraction__169 != result_fraction__871;
  assign eq_160082 = x_bexp__459 == high_exp__282;
  assign eq_160083 = x_fraction__459 == result_fraction__685;
  assign eq_160084 = prod_bexp__227 == high_exp__283;
  assign eq_160085 = prod_fraction__169 == result_fraction__686;
  assign result_exp__193 = exp__269[8:0];
  assign result_exp__34 = result_exp__33 & {9{$signed(exp__47) > $signed(10'h000)}};
  assign high_exp__153 = 8'hff;
  assign result_fraction__556 = 23'h00_0000;
  assign result_fraction__555 = 23'h00_0000;
  assign result_exp__75 = result_exp__73 & {9{$signed(exp__105) > $signed(10'h000)}};
  assign result_exp__135 = result_exp__133 & {9{$signed(exp__187) > $signed(10'h000)}};
  assign high_exp__287 = 8'hff;
  assign result_fraction__690 = 23'h00_0000;
  assign result_fraction__689 = 23'h00_0000;
  assign result_exp__195 = result_exp__193 & {9{$signed(exp__269) > $signed(10'h000)}};
  assign high_exp__86 = 8'hff;
  assign result_fraction__756 = 23'h00_0000;
  assign high_exp__87 = 8'hff;
  assign result_fraction__757 = 23'h00_0000;
  assign result_fraction__488 = 23'h00_0000;
  assign result_fraction__489 = 23'h00_0000;
  assign wide_exponent__32 = wide_exponent__31[8:0] & {9{~wide_exponent__31[9]}};
  assign has_pos_inf__10 = ~(x_bexp__86 != high_exp__365 | ne_160043 | x_sign__22) | ~(prod_bexp__42 != high_exp__366 | ne_160045 | prod_sign__10);
  assign has_neg_inf__10 = eq_160046 & eq_160047 & x_sign__22 | eq_160048 & eq_160049 & prod_sign__10;
  assign high_exp__150 = 8'hff;
  assign result_fraction__789 = 23'h00_0000;
  assign high_exp__151 = 8'hff;
  assign result_fraction__790 = 23'h00_0000;
  assign result_fraction__553 = 23'h00_0000;
  assign result_fraction__554 = 23'h00_0000;
  assign wide_exponent__68 = wide_exponent__66[8:0] & {9{~wide_exponent__66[9]}};
  assign has_pos_inf__22 = ~(x_bexp__171 != high_exp__397 | ne_160055 | x_sign__43) | ~(prod_bexp__83 != high_exp__398 | ne_160057 | prod_sign__21);
  assign has_neg_inf__22 = eq_160058 & eq_160059 & x_sign__43 | eq_160060 & eq_160061 & prod_sign__21;
  assign eq_160149 = x_bexp__173 == high_exp__153;
  assign ne_160150 = x_fraction__173 != result_fraction__556;
  assign high_exp__215 = 8'hff;
  assign result_fraction__822 = 23'h00_0000;
  assign high_exp__216 = 8'hff;
  assign result_fraction__823 = 23'h00_0000;
  assign result_fraction__618 = 23'h00_0000;
  assign result_fraction__619 = 23'h00_0000;
  assign wide_exponent__125 = wide_exponent__123[8:0] & {9{~wide_exponent__123[9]}};
  assign has_pos_inf__41 = ~(x_bexp__315 != high_exp__429 | ne_160067 | x_sign__79) | ~(prod_bexp__155 != high_exp__430 | ne_160069 | prod_sign__39);
  assign has_neg_inf__41 = eq_160070 & eq_160071 & x_sign__79 | eq_160072 & eq_160073 & prod_sign__39;
  assign high_exp__284 = 8'hff;
  assign result_fraction__855 = 23'h00_0000;
  assign high_exp__285 = 8'hff;
  assign result_fraction__856 = 23'h00_0000;
  assign result_fraction__687 = 23'h00_0000;
  assign result_fraction__688 = 23'h00_0000;
  assign wide_exponent__182 = wide_exponent__180[8:0] & {9{~wide_exponent__180[9]}};
  assign has_pos_inf__60 = ~(x_bexp__459 != high_exp__461 | ne_160079 | x_sign__115) | ~(prod_bexp__227 != high_exp__462 | ne_160081 | prod_sign__57);
  assign has_neg_inf__60 = eq_160082 & eq_160083 & x_sign__115 | eq_160084 & eq_160085 & prod_sign__57;
  assign is_result_nan__60 = x_bexp__461 == high_exp__287;
  assign ne_160177 = x_fraction__461 != result_fraction__690;
  assign wide_exponent__6 = wide_exponent__5[8:0] & {9{~wide_exponent__5[9]}};
  assign eq_160181 = x_bexp__14 == high_exp__86;
  assign ne_160182 = x_fraction__14 != result_fraction__756;
  assign eq_160183 = prod_bexp__6 == high_exp__87;
  assign ne_160184 = prod_fraction__4 != result_fraction__757;
  assign and_reduce_160195 = &result_exp__34[7:0];
  assign wide_exponent__69 = wide_exponent__67[8:0] & {9{~wide_exponent__67[9]}};
  assign eq_160197 = x_bexp__172 == high_exp__150;
  assign ne_160198 = x_fraction__172 != result_fraction__789;
  assign eq_160199 = prod_bexp__84 == high_exp__151;
  assign ne_160200 = prod_fraction__62 != result_fraction__790;
  assign is_result_nan__48 = eq_160149 & ne_160150;
  assign has_inf_arg__25 = eq_160149 & x_fraction__173 == result_fraction__555;
  assign and_reduce_160213 = &result_exp__75[7:0];
  assign wide_exponent__126 = wide_exponent__124[8:0] & {9{~wide_exponent__124[9]}};
  assign eq_160215 = x_bexp__316 == high_exp__215;
  assign ne_160216 = x_fraction__316 != result_fraction__822;
  assign eq_160217 = prod_bexp__156 == high_exp__216;
  assign ne_160218 = prod_fraction__116 != result_fraction__823;
  assign and_reduce_160229 = &result_exp__135[7:0];
  assign wide_exponent__183 = wide_exponent__181[8:0] & {9{~wide_exponent__181[9]}};
  assign eq_160231 = x_bexp__460 == high_exp__284;
  assign ne_160232 = x_fraction__460 != result_fraction__855;
  assign eq_160233 = prod_bexp__228 == high_exp__285;
  assign ne_160234 = prod_fraction__170 != result_fraction__856;
  assign is_result_nan__126 = is_result_nan__60 & ne_160177;
  assign has_inf_arg__65 = is_result_nan__60 & x_fraction__461 == result_fraction__689;
  assign and_reduce_160247 = &result_exp__195[7:0];
  assign is_result_nan__21 = eq_160046 & ne_160043 | eq_160048 & ne_160045 | has_pos_inf__10 & has_neg_inf__10;
  assign is_operand_inf__10 = eq_160046 & eq_160047 | eq_160048 & eq_160049;
  assign and_reduce_160260 = &wide_exponent__32[7:0];
  assign high_exp__90 = 8'hff;
  assign is_result_nan__46 = eq_160058 & ne_160055 | eq_160060 & ne_160057 | has_pos_inf__22 & has_neg_inf__22;
  assign is_operand_inf__22 = eq_160058 & eq_160059 | eq_160060 & eq_160061;
  assign and_reduce_160275 = &wide_exponent__68[7:0];
  assign high_exp__155 = 8'hff;
  assign is_result_nan__85 = eq_160070 & ne_160067 | eq_160072 & ne_160069 | has_pos_inf__41 & has_neg_inf__41;
  assign is_operand_inf__41 = eq_160070 & eq_160071 | eq_160072 & eq_160073;
  assign and_reduce_160290 = &wide_exponent__125[7:0];
  assign high_exp__219 = 8'hff;
  assign is_result_nan__124 = eq_160082 & ne_160079 | eq_160084 & ne_160081 | has_pos_inf__60 & has_neg_inf__60;
  assign is_operand_inf__60 = eq_160082 & eq_160083 | eq_160084 & eq_160085;
  assign and_reduce_160305 = &wide_exponent__182[7:0];
  assign high_exp__289 = 8'hff;
  assign is_result_nan__4 = eq_160181 & ne_160182 | eq_160183 & ne_160184;
  assign is_operand_inf__2 = eq_160181 & x_fraction__14 == result_fraction__488 | eq_160183 & prod_fraction__4 == result_fraction__489;
  assign and_reduce_160313 = &wide_exponent__6[7:0];
  assign fraction_shift__368 = 3'h3;
  assign fraction_shift__231 = 3'h4;
  assign is_subnormal__11 = $signed(exp__47) <= $signed(10'h000);
  assign high_exp__88 = 8'hff;
  assign result_exp__35 = is_result_nan__44 | has_inf_arg__24 | result_exp__34[8] | and_reduce_160195 ? high_exp__90 : result_exp__34[7:0];
  assign is_result_nan__47 = eq_160197 & ne_160198 | eq_160199 & ne_160200;
  assign is_operand_inf__23 = eq_160197 & x_fraction__172 == result_fraction__553 | eq_160199 & prod_fraction__62 == result_fraction__554;
  assign and_reduce_160326 = &wide_exponent__69[7:0];
  assign fraction_shift__386 = 3'h3;
  assign fraction_shift__266 = 3'h4;
  assign is_subnormal__25 = $signed(exp__105) <= $signed(10'h000);
  assign high_exp__152 = 8'hff;
  assign result_exp__77 = is_result_nan__48 | has_inf_arg__25 | result_exp__75[8] | and_reduce_160213 ? high_exp__155 : result_exp__75[7:0];
  assign is_result_nan__86 = eq_160215 & ne_160216 | eq_160217 & ne_160218;
  assign is_operand_inf__42 = eq_160215 & x_fraction__316 == result_fraction__618 | eq_160217 & prod_fraction__116 == result_fraction__619;
  assign and_reduce_160339 = &wide_exponent__126[7:0];
  assign fraction_shift__404 = 3'h3;
  assign fraction_shift__301 = 3'h4;
  assign is_subnormal__45 = $signed(exp__187) <= $signed(10'h000);
  assign high_exp__217 = 8'hff;
  assign result_exp__137 = is_result_nan__122 | has_inf_arg__64 | result_exp__135[8] | and_reduce_160229 ? high_exp__219 : result_exp__135[7:0];
  assign is_result_nan__125 = eq_160231 & ne_160232 | eq_160233 & ne_160234;
  assign is_operand_inf__61 = eq_160231 & x_fraction__460 == result_fraction__687 | eq_160233 & prod_fraction__170 == result_fraction__688;
  assign and_reduce_160352 = &wide_exponent__183[7:0];
  assign fraction_shift__422 = 3'h3;
  assign fraction_shift__336 = 3'h4;
  assign is_subnormal__65 = $signed(exp__269) <= $signed(10'h000);
  assign high_exp__286 = 8'hff;
  assign result_exp__197 = is_result_nan__126 | has_inf_arg__65 | result_exp__195[8] | and_reduce_160247 ? high_exp__289 : result_exp__195[7:0];
  assign fraction_shift__369 = 3'h3;
  assign fraction_shift__232 = 3'h4;
  assign high_exp__89 = 8'hff;
  assign fraction_shift__33 = rounding_carry__10 ? fraction_shift__231 : fraction_shift__368;
  assign result_sign__403 = 1'h0;
  assign result_exponent__11 = is_result_nan__21 | is_operand_inf__10 | wide_exponent__32[8] | and_reduce_160260 ? high_exp__88 : wide_exponent__32[7:0];
  assign result_sign__404 = 1'h0;
  assign fraction_shift__387 = 3'h3;
  assign fraction_shift__267 = 3'h4;
  assign high_exp__154 = 8'hff;
  assign fraction_shift__68 = rounding_carry__22 ? fraction_shift__266 : fraction_shift__386;
  assign result_sign__500 = 1'h0;
  assign result_exponent__22 = is_result_nan__46 | is_operand_inf__22 | wide_exponent__68[8] | and_reduce_160275 ? high_exp__152 : wide_exponent__68[7:0];
  assign result_sign__501 = 1'h0;
  assign fraction_shift__405 = 3'h3;
  assign fraction_shift__302 = 3'h4;
  assign high_exp__218 = 8'hff;
  assign fraction_shift__125 = rounding_carry__41 ? fraction_shift__301 : fraction_shift__404;
  assign result_sign__593 = 1'h0;
  assign result_exponent__41 = is_result_nan__85 | is_operand_inf__41 | wide_exponent__125[8] | and_reduce_160290 ? high_exp__217 : wide_exponent__125[7:0];
  assign result_sign__594 = 1'h0;
  assign fraction_shift__423 = 3'h3;
  assign fraction_shift__337 = 3'h4;
  assign high_exp__288 = 8'hff;
  assign fraction_shift__182 = rounding_carry__60 ? fraction_shift__336 : fraction_shift__422;
  assign result_sign__699 = 1'h0;
  assign result_exponent__60 = is_result_nan__124 | is_operand_inf__60 | wide_exponent__182[8] | and_reduce_160305 ? high_exp__286 : wide_exponent__182[7:0];
  assign result_sign__700 = 1'h0;
  assign fraction_shift__6 = rounding_carry__2 ? fraction_shift__232 : fraction_shift__369;
  assign result_sign__405 = 1'h0;
  assign result_exponent__1 = is_result_nan__4 | is_operand_inf__2 | wide_exponent__6[8] | and_reduce_160313 ? high_exp__89 : wide_exponent__6[7:0];
  assign shrl_160412 = rounded_fraction__10 >> fraction_shift__33;
  assign concat_160416 = {result_sign__404, ~result_exp__35};
  assign fraction_shift__69 = rounding_carry__23 ? fraction_shift__267 : fraction_shift__387;
  assign result_sign__502 = 1'h0;
  assign result_exponent__23 = is_result_nan__47 | is_operand_inf__23 | wide_exponent__69[8] | and_reduce_160326 ? high_exp__154 : wide_exponent__69[7:0];
  assign shrl_160421 = rounded_fraction__22 >> fraction_shift__68;
  assign concat_160425 = {result_sign__501, ~result_exp__77};
  assign fraction_shift__126 = rounding_carry__42 ? fraction_shift__302 : fraction_shift__405;
  assign result_sign__595 = 1'h0;
  assign result_exponent__42 = is_result_nan__86 | is_operand_inf__42 | wide_exponent__126[8] | and_reduce_160339 ? high_exp__218 : wide_exponent__126[7:0];
  assign shrl_160430 = rounded_fraction__41 >> fraction_shift__125;
  assign concat_160434 = {result_sign__594, ~result_exp__137};
  assign fraction_shift__183 = rounding_carry__61 ? fraction_shift__337 : fraction_shift__423;
  assign result_sign__701 = 1'h0;
  assign result_exponent__61 = is_result_nan__125 | is_operand_inf__61 | wide_exponent__183[8] | and_reduce_160352 ? high_exp__288 : wide_exponent__183[7:0];
  assign shrl_160439 = rounded_fraction__60 >> fraction_shift__182;
  assign concat_160443 = {result_sign__700, ~result_exp__197};
  assign shrl_160444 = rounded_fraction__2 >> fraction_shift__6;
  assign result_fraction__63 = shrl_160412[22:0];
  assign result_fraction__66 = fraction__106[22:0];
  assign sum__11 = {result_sign__403, result_exponent__11} + concat_160416;
  assign shrl_160452 = rounded_fraction__23 >> fraction_shift__69;
  assign result_fraction__136 = shrl_160421[22:0];
  assign result_fraction__142 = fraction__230[22:0];
  assign sum__24 = {result_sign__500, result_exponent__22} + concat_160425;
  assign shrl_160460 = rounded_fraction__42 >> fraction_shift__126;
  assign result_fraction__253 = shrl_160430[22:0];
  assign result_fraction__259 = fraction__409[22:0];
  assign sum__43 = {result_sign__593, result_exponent__41} + concat_160434;
  assign shrl_160468 = rounded_fraction__61 >> fraction_shift__183;
  assign result_fraction__370 = shrl_160439[22:0];
  assign result_fraction__376 = fraction__588[22:0];
  assign sum__62 = {result_sign__699, result_exponent__60} + concat_160443;
  assign result_fraction__10 = shrl_160444[22:0];
  assign sum__3 = {result_sign__405, result_exponent__1} + concat_160416;
  assign result_fraction__64 = result_fraction__63 & {23{~(is_operand_inf__10 | wide_exponent__32[8] | and_reduce_160260 | ~((|wide_exponent__32[8:1]) | wide_exponent__32[0]))}};
  assign nan_fraction__83 = 23'h40_0000;
  assign result_fraction__67 = result_fraction__66 & {23{~(has_inf_arg__24 | result_exp__34[8] | and_reduce_160195 | is_subnormal__11)}};
  assign nan_fraction__85 = 23'h40_0000;
  assign result_fraction__137 = shrl_160452[22:0];
  assign sum__25 = {result_sign__502, result_exponent__23} + concat_160425;
  assign result_fraction__138 = result_fraction__136 & {23{~(is_operand_inf__22 | wide_exponent__68[8] | and_reduce_160275 | ~((|wide_exponent__68[8:1]) | wide_exponent__68[0]))}};
  assign nan_fraction__110 = 23'h40_0000;
  assign result_fraction__144 = result_fraction__142 & {23{~(has_inf_arg__25 | result_exp__75[8] | and_reduce_160213 | is_subnormal__25)}};
  assign nan_fraction__112 = 23'h40_0000;
  assign result_fraction__254 = shrl_160460[22:0];
  assign sum__44 = {result_sign__595, result_exponent__42} + concat_160434;
  assign result_fraction__255 = result_fraction__253 & {23{~(is_operand_inf__41 | wide_exponent__125[8] | and_reduce_160290 | ~((|wide_exponent__125[8:1]) | wide_exponent__125[0]))}};
  assign nan_fraction__137 = 23'h40_0000;
  assign result_fraction__261 = result_fraction__259 & {23{~(has_inf_arg__64 | result_exp__135[8] | and_reduce_160229 | is_subnormal__45)}};
  assign nan_fraction__139 = 23'h40_0000;
  assign result_fraction__371 = shrl_160468[22:0];
  assign sum__63 = {result_sign__701, result_exponent__61} + concat_160443;
  assign result_fraction__372 = result_fraction__370 & {23{~(is_operand_inf__60 | wide_exponent__182[8] | and_reduce_160305 | ~((|wide_exponent__182[8:1]) | wide_exponent__182[0]))}};
  assign nan_fraction__166 = 23'h40_0000;
  assign result_fraction__378 = result_fraction__376 & {23{~(has_inf_arg__65 | result_exp__195[8] | and_reduce_160247 | is_subnormal__65)}};
  assign nan_fraction__168 = 23'h40_0000;
  assign result_fraction__11 = result_fraction__10 & {23{~(is_operand_inf__2 | wide_exponent__6[8] | and_reduce_160313 | ~((|wide_exponent__6[8:1]) | wide_exponent__6[0]))}};
  assign nan_fraction__84 = 23'h40_0000;
  assign result_fraction__65 = is_result_nan__21 ? nan_fraction__83 : result_fraction__64;
  assign result_fraction__68 = is_result_nan__44 ? nan_fraction__85 : result_fraction__67;
  assign prod_bexp__46 = sum__11[8] ? result_exp__35 : result_exponent__11;
  assign x_bexp__692 = 8'h00;
  assign result_fraction__139 = result_fraction__137 & {23{~(is_operand_inf__23 | wide_exponent__69[8] | and_reduce_160326 | ~((|wide_exponent__69[8:1]) | wide_exponent__69[0]))}};
  assign nan_fraction__111 = 23'h40_0000;
  assign result_fraction__140 = is_result_nan__46 ? nan_fraction__110 : result_fraction__138;
  assign result_fraction__146 = is_result_nan__48 ? nan_fraction__112 : result_fraction__144;
  assign prod_bexp__91 = sum__24[8] ? result_exp__77 : result_exponent__22;
  assign x_bexp__693 = 8'h00;
  assign result_fraction__256 = result_fraction__254 & {23{~(is_operand_inf__42 | wide_exponent__126[8] | and_reduce_160339 | ~((|wide_exponent__126[8:1]) | wide_exponent__126[0]))}};
  assign nan_fraction__138 = 23'h40_0000;
  assign result_fraction__257 = is_result_nan__85 ? nan_fraction__137 : result_fraction__255;
  assign result_fraction__263 = is_result_nan__122 ? nan_fraction__139 : result_fraction__261;
  assign prod_bexp__163 = sum__43[8] ? result_exp__137 : result_exponent__41;
  assign x_bexp__694 = 8'h00;
  assign result_fraction__373 = result_fraction__371 & {23{~(is_operand_inf__61 | wide_exponent__183[8] | and_reduce_160352 | ~((|wide_exponent__183[8:1]) | wide_exponent__183[0]))}};
  assign nan_fraction__167 = 23'h40_0000;
  assign result_fraction__374 = is_result_nan__124 ? nan_fraction__166 : result_fraction__372;
  assign result_fraction__380 = is_result_nan__126 ? nan_fraction__168 : result_fraction__378;
  assign prod_bexp__235 = sum__62[8] ? result_exp__197 : result_exponent__60;
  assign x_bexp__695 = 8'h00;
  assign high_exp__351 = 8'hff;
  assign high_exp__352 = 8'hff;
  assign result_fraction__12 = is_result_nan__4 ? nan_fraction__84 : result_fraction__11;
  assign prod_bexp__10 = sum__3[8] ? result_exp__35 : result_exponent__1;
  assign x_bexp__696 = 8'h00;
  assign fraction_is_zero__10 = add_159320 == 26'h000_0000 & xddend_y__10[2:0] == 3'h0;
  assign prod_fraction__33 = sum__11[8] ? result_fraction__68 : result_fraction__65;
  assign incremented_sum__80 = sum__11[7:0] + 8'h01;
  assign high_exp__383 = 8'hff;
  assign high_exp__384 = 8'hff;
  assign result_fraction__141 = is_result_nan__47 ? nan_fraction__111 : result_fraction__139;
  assign prod_bexp__92 = sum__25[8] ? result_exp__77 : result_exponent__23;
  assign x_bexp__697 = 8'h00;
  assign fraction_is_zero__22 = add_159323 == 26'h000_0000 & xddend_y__21[2:0] == 3'h0;
  assign prod_fraction__67 = sum__24[8] ? result_fraction__146 : result_fraction__140;
  assign incremented_sum__98 = sum__24[7:0] + 8'h01;
  assign high_exp__415 = 8'hff;
  assign high_exp__416 = 8'hff;
  assign result_fraction__258 = is_result_nan__86 ? nan_fraction__138 : result_fraction__256;
  assign prod_bexp__164 = sum__44[8] ? result_exp__137 : result_exponent__42;
  assign x_bexp__698 = 8'h00;
  assign fraction_is_zero__41 = add_159326 == 26'h000_0000 & xddend_y__39[2:0] == 3'h0;
  assign prod_fraction__121 = sum__43[8] ? result_fraction__263 : result_fraction__257;
  assign incremented_sum__116 = sum__43[7:0] + 8'h01;
  assign high_exp__447 = 8'hff;
  assign high_exp__448 = 8'hff;
  assign result_fraction__375 = is_result_nan__125 ? nan_fraction__167 : result_fraction__373;
  assign prod_bexp__236 = sum__63[8] ? result_exp__197 : result_exponent__61;
  assign x_bexp__699 = 8'h00;
  assign fraction_is_zero__60 = add_159329 == 26'h000_0000 & xddend_y__57[2:0] == 3'h0;
  assign prod_fraction__175 = sum__62[8] ? result_fraction__380 : result_fraction__374;
  assign incremented_sum__134 = sum__62[7:0] + 8'h01;
  assign fraction_is_zero__2 = add_159330 == 26'h000_0000 & xddend_y__2[2:0] == 3'h0;
  assign prod_fraction__7 = sum__3[8] ? result_fraction__68 : result_fraction__12;
  assign incremented_sum__81 = sum__3[7:0] + 8'h01;
  assign wide_y__22 = {2'h1, prod_fraction__33, 3'h0};
  assign x_bexpbs_difference__12 = sum__11[8] ? incremented_sum__80 : ~sum__11[7:0];
  assign fraction_is_zero__23 = add_159333 == 26'h000_0000 & xddend_y__22[2:0] == 3'h0;
  assign prod_fraction__68 = sum__25[8] ? result_fraction__146 : result_fraction__141;
  assign incremented_sum__99 = sum__25[7:0] + 8'h01;
  assign wide_y__47 = {2'h1, prod_fraction__67, 3'h0};
  assign x_bexpbs_difference__23 = sum__24[8] ? incremented_sum__98 : ~sum__24[7:0];
  assign fraction_is_zero__42 = add_159336 == 26'h000_0000 & xddend_y__40[2:0] == 3'h0;
  assign prod_fraction__122 = sum__44[8] ? result_fraction__263 : result_fraction__258;
  assign incremented_sum__117 = sum__44[7:0] + 8'h01;
  assign wide_y__85 = {2'h1, prod_fraction__121, 3'h0};
  assign x_bexpbs_difference__41 = sum__43[8] ? incremented_sum__116 : ~sum__43[7:0];
  assign fraction_is_zero__61 = add_159339 == 26'h000_0000 & xddend_y__58[2:0] == 3'h0;
  assign prod_fraction__176 = sum__63[8] ? result_fraction__380 : result_fraction__375;
  assign incremented_sum__135 = sum__63[7:0] + 8'h01;
  assign wide_y__123 = {2'h1, prod_fraction__175, 3'h0};
  assign x_bexpbs_difference__59 = sum__62[8] ? incremented_sum__134 : ~sum__62[7:0];
  assign wide_y__5 = {2'h1, prod_fraction__7, 3'h0};
  assign x_bexpbs_difference__3 = sum__3[8] ? incremented_sum__81 : ~sum__3[7:0];
  assign concat_160695 = {~(add_159320[25] | fraction_is_zero__10), add_159320[25], fraction_is_zero__10};
  assign x_bexp__94 = sum__11[8] ? result_exponent__11 : result_exp__35;
  assign x_bexp__700 = 8'h00;
  assign wide_y__23 = wide_y__22 & {28{prod_bexp__46 != x_bexp__692}};
  assign sub_160701 = 8'h1c - x_bexpbs_difference__12;
  assign wide_y__48 = {2'h1, prod_fraction__68, 3'h0};
  assign x_bexpbs_difference__24 = sum__25[8] ? incremented_sum__99 : ~sum__25[7:0];
  assign concat_160709 = {~(add_159323[25] | fraction_is_zero__22), add_159323[25], fraction_is_zero__22};
  assign x_bexp__187 = sum__24[8] ? result_exponent__22 : result_exp__77;
  assign x_bexp__701 = 8'h00;
  assign wide_y__49 = wide_y__47 & {28{prod_bexp__91 != x_bexp__693}};
  assign sub_160715 = 8'h1c - x_bexpbs_difference__23;
  assign wide_y__86 = {2'h1, prod_fraction__122, 3'h0};
  assign x_bexpbs_difference__42 = sum__44[8] ? incremented_sum__117 : ~sum__44[7:0];
  assign concat_160723 = {~(add_159326[25] | fraction_is_zero__41), add_159326[25], fraction_is_zero__41};
  assign x_bexp__331 = sum__43[8] ? result_exponent__41 : result_exp__137;
  assign x_bexp__702 = 8'h00;
  assign wide_y__87 = wide_y__85 & {28{prod_bexp__163 != x_bexp__694}};
  assign sub_160729 = 8'h1c - x_bexpbs_difference__41;
  assign wide_y__124 = {2'h1, prod_fraction__176, 3'h0};
  assign x_bexpbs_difference__60 = sum__63[8] ? incremented_sum__135 : ~sum__63[7:0];
  assign concat_160737 = {~(add_159329[25] | fraction_is_zero__60), add_159329[25], fraction_is_zero__60};
  assign x_bexp__475 = sum__62[8] ? result_exponent__60 : result_exp__197;
  assign x_bexp__703 = 8'h00;
  assign wide_y__125 = wide_y__123 & {28{prod_bexp__235 != x_bexp__695}};
  assign sub_160743 = 8'h1c - x_bexpbs_difference__59;
  assign concat_160744 = {~(add_159330[25] | fraction_is_zero__2), add_159330[25], fraction_is_zero__2};
  assign has_pos_inf__2 = ~(x_bexp__14 != high_exp__351 | ne_160182 | x_sign__4) | ~(prod_bexp__6 != high_exp__352 | ne_160184 | prod_sign__2);
  assign x_bexp__22 = sum__3[8] ? result_exponent__1 : result_exp__35;
  assign x_bexp__704 = 8'h00;
  assign wide_y__6 = wide_y__5 & {28{prod_bexp__10 != x_bexp__696}};
  assign sub_160751 = 8'h1c - x_bexpbs_difference__3;
  assign result_sign__52 = x_sign__22 & prod_sign__10 & concat_160695[0] | ~prod_sign__10 & concat_160695[1] | prod_sign__10 & concat_160695[2];
  assign x_fraction__94 = sum__11[8] ? result_fraction__65 : result_fraction__68;
  assign dropped__11 = sub_160701 >= 8'h1c ? 28'h000_0000 : wide_y__23 << sub_160701;
  assign concat_160759 = {~(add_159333[25] | fraction_is_zero__23), add_159333[25], fraction_is_zero__23};
  assign has_pos_inf__23 = ~(x_bexp__172 != high_exp__383 | ne_160198 | x_sign__44) | ~(prod_bexp__84 != high_exp__384 | ne_160200 | prod_sign__22);
  assign x_bexp__188 = sum__25[8] ? result_exponent__23 : result_exp__77;
  assign x_bexp__705 = 8'h00;
  assign wide_y__50 = wide_y__48 & {28{prod_bexp__92 != x_bexp__697}};
  assign sub_160766 = 8'h1c - x_bexpbs_difference__24;
  assign x_sign__45 = array_index_159490[31:31];
  assign result_sign__112 = x_sign__43 & prod_sign__21 & concat_160709[0] | ~prod_sign__21 & concat_160709[1] | prod_sign__21 & concat_160709[2];
  assign x_fraction__187 = sum__24[8] ? result_fraction__140 : result_fraction__146;
  assign dropped__24 = sub_160715 >= 8'h1c ? 28'h000_0000 : wide_y__49 << sub_160715;
  assign concat_160775 = {~(add_159336[25] | fraction_is_zero__42), add_159336[25], fraction_is_zero__42};
  assign has_pos_inf__42 = ~(x_bexp__316 != high_exp__415 | ne_160216 | x_sign__80) | ~(prod_bexp__156 != high_exp__416 | ne_160218 | prod_sign__40);
  assign x_bexp__332 = sum__44[8] ? result_exponent__42 : result_exp__137;
  assign x_bexp__706 = 8'h00;
  assign wide_y__88 = wide_y__86 & {28{prod_bexp__164 != x_bexp__698}};
  assign sub_160782 = 8'h1c - x_bexpbs_difference__42;
  assign result_sign__209 = x_sign__79 & prod_sign__39 & concat_160723[0] | ~prod_sign__39 & concat_160723[1] | prod_sign__39 & concat_160723[2];
  assign x_fraction__331 = sum__43[8] ? result_fraction__257 : result_fraction__263;
  assign dropped__43 = sub_160729 >= 8'h1c ? 28'h000_0000 : wide_y__87 << sub_160729;
  assign concat_160790 = {~(add_159339[25] | fraction_is_zero__61), add_159339[25], fraction_is_zero__61};
  assign has_pos_inf__61 = ~(x_bexp__460 != high_exp__447 | ne_160232 | x_sign__116) | ~(prod_bexp__228 != high_exp__448 | ne_160234 | prod_sign__58);
  assign x_bexp__476 = sum__63[8] ? result_exponent__61 : result_exp__197;
  assign x_bexp__707 = 8'h00;
  assign wide_y__126 = wide_y__124 & {28{prod_bexp__236 != x_bexp__699}};
  assign sub_160797 = 8'h1c - x_bexpbs_difference__60;
  assign x_sign__117 = array_index_159517[31:31];
  assign result_sign__306 = x_sign__115 & prod_sign__57 & concat_160737[0] | ~prod_sign__57 & concat_160737[1] | prod_sign__57 & concat_160737[2];
  assign x_fraction__475 = sum__62[8] ? result_fraction__374 : result_fraction__380;
  assign dropped__62 = sub_160743 >= 8'h1c ? 28'h000_0000 : wide_y__125 << sub_160743;
  assign result_sign__8 = x_sign__4 & prod_sign__2 & concat_160744[0] | ~prod_sign__2 & concat_160744[1] | prod_sign__2 & concat_160744[2];
  assign x_fraction__22 = sum__3[8] ? result_fraction__12 : result_fraction__68;
  assign dropped__3 = sub_160751 >= 8'h1c ? 28'h000_0000 : wide_y__6 << sub_160751;
  assign result_sign__53 = is_operand_inf__10 ? ~has_pos_inf__10 : result_sign__52;
  assign wide_x__22 = {2'h1, x_fraction__94, 3'h0};
  assign result_sign__113 = x_sign__44 & prod_sign__22 & concat_160759[0] | ~prod_sign__22 & concat_160759[1] | prod_sign__22 & concat_160759[2];
  assign x_fraction__188 = sum__25[8] ? result_fraction__141 : result_fraction__146;
  assign dropped__25 = sub_160766 >= 8'h1c ? 28'h000_0000 : wide_y__50 << sub_160766;
  assign nand_160826 = ~(eq_160149 & ne_160150);
  assign result_sign__118 = ~x_sign__45;
  assign result_sign__114 = is_operand_inf__22 ? ~has_pos_inf__22 : result_sign__112;
  assign wide_x__47 = {2'h1, x_fraction__187, 3'h0};
  assign result_sign__210 = x_sign__80 & prod_sign__40 & concat_160775[0] | ~prod_sign__40 & concat_160775[1] | prod_sign__40 & concat_160775[2];
  assign x_fraction__332 = sum__44[8] ? result_fraction__258 : result_fraction__263;
  assign dropped__44 = sub_160782 >= 8'h1c ? 28'h000_0000 : wide_y__88 << sub_160782;
  assign result_sign__211 = is_operand_inf__41 ? ~has_pos_inf__41 : result_sign__209;
  assign wide_x__85 = {2'h1, x_fraction__331, 3'h0};
  assign result_sign__307 = x_sign__116 & prod_sign__58 & concat_160790[0] | ~prod_sign__58 & concat_160790[1] | prod_sign__58 & concat_160790[2];
  assign x_fraction__476 = sum__63[8] ? result_fraction__375 : result_fraction__380;
  assign dropped__63 = sub_160797 >= 8'h1c ? 28'h000_0000 : wide_y__126 << sub_160797;
  assign nand_160854 = ~(is_result_nan__60 & ne_160177);
  assign result_sign__312 = ~x_sign__117;
  assign result_sign__308 = is_operand_inf__60 ? ~has_pos_inf__60 : result_sign__306;
  assign wide_x__123 = {2'h1, x_fraction__475, 3'h0};
  assign result_sign__9 = is_operand_inf__2 ? ~has_pos_inf__2 : result_sign__8;
  assign wide_x__5 = {2'h1, x_fraction__22, 3'h0};
  assign result_sign__54 = ~is_result_nan__21 & result_sign__53;
  assign wide_x__23 = wide_x__22 & {28{x_bexp__94 != x_bexp__700}};
  assign result_sign__115 = is_operand_inf__23 ? ~has_pos_inf__23 : result_sign__113;
  assign wide_x__48 = {2'h1, x_fraction__188, 3'h0};
  assign result_sign__120 = nand_160826 & result_sign__118;
  assign result_sign__116 = ~is_result_nan__46 & result_sign__114;
  assign wide_x__49 = wide_x__47 & {28{x_bexp__187 != x_bexp__701}};
  assign result_sign__212 = is_operand_inf__42 ? ~has_pos_inf__42 : result_sign__210;
  assign wide_x__86 = {2'h1, x_fraction__332, 3'h0};
  assign result_sign__213 = ~is_result_nan__85 & result_sign__211;
  assign wide_x__87 = wide_x__85 & {28{x_bexp__331 != x_bexp__702}};
  assign result_sign__309 = is_operand_inf__61 ? ~has_pos_inf__61 : result_sign__307;
  assign wide_x__124 = {2'h1, x_fraction__476, 3'h0};
  assign result_sign__314 = nand_160854 & result_sign__312;
  assign result_sign__310 = ~is_result_nan__124 & result_sign__308;
  assign wide_x__125 = wide_x__123 & {28{x_bexp__475 != x_bexp__703}};
  assign result_sign__12 = nand_159126 & x_sign__41;
  assign result_sign__10 = ~is_result_nan__4 & result_sign__9;
  assign wide_x__6 = wide_x__5 & {28{x_bexp__22 != x_bexp__704}};
  assign x_sign__24 = sum__11[8] ? result_sign__54 : result_sign__110;
  assign prod_sign__11 = sum__11[8] ? result_sign__110 : result_sign__54;
  assign neg_160911 = -wide_x__23;
  assign sticky__35 = {27'h000_0000, dropped__11[27:3] != 25'h000_0000};
  assign result_sign__121 = nand_160826 & x_sign__45;
  assign result_sign__117 = ~is_result_nan__47 & result_sign__115;
  assign wide_x__50 = wide_x__48 & {28{x_bexp__188 != x_bexp__705}};
  assign x_sign__47 = sum__24[8] ? result_sign__116 : result_sign__120;
  assign prod_sign__23 = sum__24[8] ? result_sign__120 : result_sign__116;
  assign neg_160921 = -wide_x__49;
  assign sticky__76 = {27'h000_0000, dropped__24[27:3] != 25'h000_0000};
  assign result_sign__218 = nand_159152 & x_sign__113;
  assign result_sign__214 = ~is_result_nan__86 & result_sign__212;
  assign wide_x__88 = wide_x__86 & {28{x_bexp__332 != x_bexp__706}};
  assign x_sign__83 = sum__43[8] ? result_sign__213 : result_sign__304;
  assign prod_sign__41 = sum__43[8] ? result_sign__304 : result_sign__213;
  assign neg_160931 = -wide_x__87;
  assign sticky__135 = {27'h000_0000, dropped__43[27:3] != 25'h000_0000};
  assign result_sign__315 = nand_160854 & x_sign__117;
  assign result_sign__311 = ~is_result_nan__125 & result_sign__309;
  assign wide_x__126 = wide_x__124 & {28{x_bexp__476 != x_bexp__707}};
  assign x_sign__119 = sum__62[8] ? result_sign__310 : result_sign__314;
  assign prod_sign__59 = sum__62[8] ? result_sign__314 : result_sign__310;
  assign neg_160941 = -wide_x__125;
  assign sticky__194 = {27'h000_0000, dropped__62[27:3] != 25'h000_0000};
  assign x_sign__6 = sum__3[8] ? result_sign__10 : result_sign__12;
  assign prod_sign__3 = sum__3[8] ? result_sign__12 : result_sign__10;
  assign neg_160946 = -wide_x__6;
  assign sticky__9 = {27'h000_0000, dropped__3[27:3] != 25'h000_0000};
  assign xddend_y__11 = (x_bexpbs_difference__12 >= 8'h1c ? 28'h000_0000 : wide_y__23 >> x_bexpbs_difference__12) | sticky__35;
  assign x_sign__48 = sum__25[8] ? result_sign__117 : result_sign__121;
  assign prod_sign__24 = sum__25[8] ? result_sign__121 : result_sign__117;
  assign neg_160955 = -wide_x__50;
  assign sticky__77 = {27'h000_0000, dropped__25[27:3] != 25'h000_0000};
  assign xddend_y__23 = (x_bexpbs_difference__23 >= 8'h1c ? 28'h000_0000 : wide_y__49 >> x_bexpbs_difference__23) | sticky__76;
  assign x_sign__84 = sum__44[8] ? result_sign__214 : result_sign__218;
  assign prod_sign__42 = sum__44[8] ? result_sign__218 : result_sign__214;
  assign neg_160964 = -wide_x__88;
  assign sticky__136 = {27'h000_0000, dropped__44[27:3] != 25'h000_0000};
  assign xddend_y__41 = (x_bexpbs_difference__41 >= 8'h1c ? 28'h000_0000 : wide_y__87 >> x_bexpbs_difference__41) | sticky__135;
  assign x_sign__120 = sum__63[8] ? result_sign__311 : result_sign__315;
  assign prod_sign__60 = sum__63[8] ? result_sign__315 : result_sign__311;
  assign neg_160973 = -wide_x__126;
  assign sticky__195 = {27'h000_0000, dropped__63[27:3] != 25'h000_0000};
  assign xddend_y__59 = (x_bexpbs_difference__59 >= 8'h1c ? 28'h000_0000 : wide_y__125 >> x_bexpbs_difference__59) | sticky__194;
  assign xddend_y__3 = (x_bexpbs_difference__3 >= 8'h1c ? 28'h000_0000 : wide_y__6 >> x_bexpbs_difference__3) | sticky__9;
  assign sel_160984 = x_sign__24 ^ prod_sign__11 ? neg_160911[27:3] : wide_x__23[27:3];
  assign result_sign__980 = 1'h0;
  assign xddend_y__24 = (x_bexpbs_difference__24 >= 8'h1c ? 28'h000_0000 : wide_y__50 >> x_bexpbs_difference__24) | sticky__77;
  assign sel_160991 = x_sign__47 ^ prod_sign__23 ? neg_160921[27:3] : wide_x__49[27:3];
  assign result_sign__981 = 1'h0;
  assign xddend_y__42 = (x_bexpbs_difference__42 >= 8'h1c ? 28'h000_0000 : wide_y__88 >> x_bexpbs_difference__42) | sticky__136;
  assign sel_160998 = x_sign__83 ^ prod_sign__41 ? neg_160931[27:3] : wide_x__87[27:3];
  assign result_sign__982 = 1'h0;
  assign xddend_y__60 = (x_bexpbs_difference__60 >= 8'h1c ? 28'h000_0000 : wide_y__126 >> x_bexpbs_difference__60) | sticky__195;
  assign sel_161005 = x_sign__119 ^ prod_sign__59 ? neg_160941[27:3] : wide_x__125[27:3];
  assign result_sign__983 = 1'h0;
  assign sel_161008 = x_sign__6 ^ prod_sign__3 ? neg_160946[27:3] : wide_x__6[27:3];
  assign result_sign__984 = 1'h0;
  assign sel_161013 = x_sign__48 ^ prod_sign__24 ? neg_160955[27:3] : wide_x__50[27:3];
  assign result_sign__985 = 1'h0;
  assign sel_161018 = x_sign__84 ^ prod_sign__42 ? neg_160964[27:3] : wide_x__88[27:3];
  assign result_sign__986 = 1'h0;
  assign sel_161023 = x_sign__120 ^ prod_sign__60 ? neg_160973[27:3] : wide_x__126[27:3];
  assign result_sign__987 = 1'h0;
  assign add_161030 = {{1{sel_160984[24]}}, sel_160984} + {result_sign__980, xddend_y__11[27:3]};
  assign add_161033 = {{1{sel_160991[24]}}, sel_160991} + {result_sign__981, xddend_y__23[27:3]};
  assign add_161036 = {{1{sel_160998[24]}}, sel_160998} + {result_sign__982, xddend_y__41[27:3]};
  assign add_161039 = {{1{sel_161005[24]}}, sel_161005} + {result_sign__983, xddend_y__59[27:3]};
  assign add_161040 = {{1{sel_161008[24]}}, sel_161008} + {result_sign__984, xddend_y__3[27:3]};
  assign add_161043 = {{1{sel_161013[24]}}, sel_161013} + {result_sign__985, xddend_y__24[27:3]};
  assign add_161046 = {{1{sel_161018[24]}}, sel_161018} + {result_sign__986, xddend_y__42[27:3]};
  assign add_161049 = {{1{sel_161023[24]}}, sel_161023} + {result_sign__987, xddend_y__60[27:3]};
  assign concat_161054 = {add_161030[24:0], xddend_y__11[2:0]};
  assign concat_161057 = {add_161033[24:0], xddend_y__23[2:0]};
  assign concat_161060 = {add_161036[24:0], xddend_y__41[2:0]};
  assign concat_161063 = {add_161039[24:0], xddend_y__59[2:0]};
  assign concat_161064 = {add_161040[24:0], xddend_y__3[2:0]};
  assign concat_161067 = {add_161043[24:0], xddend_y__24[2:0]};
  assign concat_161070 = {add_161046[24:0], xddend_y__42[2:0]};
  assign concat_161073 = {add_161049[24:0], xddend_y__60[2:0]};
  assign xbs_fraction__11 = add_161030[25] ? -concat_161054 : concat_161054;
  assign xbs_fraction__23 = add_161033[25] ? -concat_161057 : concat_161057;
  assign xbs_fraction__41 = add_161036[25] ? -concat_161060 : concat_161060;
  assign xbs_fraction__59 = add_161039[25] ? -concat_161063 : concat_161063;
  assign xbs_fraction__3 = add_161040[25] ? -concat_161064 : concat_161064;
  assign reverse_161089 = {xbs_fraction__11[0], xbs_fraction__11[1], xbs_fraction__11[2], xbs_fraction__11[3], xbs_fraction__11[4], xbs_fraction__11[5], xbs_fraction__11[6], xbs_fraction__11[7], xbs_fraction__11[8], xbs_fraction__11[9], xbs_fraction__11[10], xbs_fraction__11[11], xbs_fraction__11[12], xbs_fraction__11[13], xbs_fraction__11[14], xbs_fraction__11[15], xbs_fraction__11[16], xbs_fraction__11[17], xbs_fraction__11[18], xbs_fraction__11[19], xbs_fraction__11[20], xbs_fraction__11[21], xbs_fraction__11[22], xbs_fraction__11[23], xbs_fraction__11[24], xbs_fraction__11[25], xbs_fraction__11[26], xbs_fraction__11[27]};
  assign xbs_fraction__24 = add_161043[25] ? -concat_161067 : concat_161067;
  assign reverse_161091 = {xbs_fraction__23[0], xbs_fraction__23[1], xbs_fraction__23[2], xbs_fraction__23[3], xbs_fraction__23[4], xbs_fraction__23[5], xbs_fraction__23[6], xbs_fraction__23[7], xbs_fraction__23[8], xbs_fraction__23[9], xbs_fraction__23[10], xbs_fraction__23[11], xbs_fraction__23[12], xbs_fraction__23[13], xbs_fraction__23[14], xbs_fraction__23[15], xbs_fraction__23[16], xbs_fraction__23[17], xbs_fraction__23[18], xbs_fraction__23[19], xbs_fraction__23[20], xbs_fraction__23[21], xbs_fraction__23[22], xbs_fraction__23[23], xbs_fraction__23[24], xbs_fraction__23[25], xbs_fraction__23[26], xbs_fraction__23[27]};
  assign xbs_fraction__42 = add_161046[25] ? -concat_161070 : concat_161070;
  assign reverse_161093 = {xbs_fraction__41[0], xbs_fraction__41[1], xbs_fraction__41[2], xbs_fraction__41[3], xbs_fraction__41[4], xbs_fraction__41[5], xbs_fraction__41[6], xbs_fraction__41[7], xbs_fraction__41[8], xbs_fraction__41[9], xbs_fraction__41[10], xbs_fraction__41[11], xbs_fraction__41[12], xbs_fraction__41[13], xbs_fraction__41[14], xbs_fraction__41[15], xbs_fraction__41[16], xbs_fraction__41[17], xbs_fraction__41[18], xbs_fraction__41[19], xbs_fraction__41[20], xbs_fraction__41[21], xbs_fraction__41[22], xbs_fraction__41[23], xbs_fraction__41[24], xbs_fraction__41[25], xbs_fraction__41[26], xbs_fraction__41[27]};
  assign xbs_fraction__60 = add_161049[25] ? -concat_161073 : concat_161073;
  assign reverse_161095 = {xbs_fraction__59[0], xbs_fraction__59[1], xbs_fraction__59[2], xbs_fraction__59[3], xbs_fraction__59[4], xbs_fraction__59[5], xbs_fraction__59[6], xbs_fraction__59[7], xbs_fraction__59[8], xbs_fraction__59[9], xbs_fraction__59[10], xbs_fraction__59[11], xbs_fraction__59[12], xbs_fraction__59[13], xbs_fraction__59[14], xbs_fraction__59[15], xbs_fraction__59[16], xbs_fraction__59[17], xbs_fraction__59[18], xbs_fraction__59[19], xbs_fraction__59[20], xbs_fraction__59[21], xbs_fraction__59[22], xbs_fraction__59[23], xbs_fraction__59[24], xbs_fraction__59[25], xbs_fraction__59[26], xbs_fraction__59[27]};
  assign reverse_161096 = {xbs_fraction__3[0], xbs_fraction__3[1], xbs_fraction__3[2], xbs_fraction__3[3], xbs_fraction__3[4], xbs_fraction__3[5], xbs_fraction__3[6], xbs_fraction__3[7], xbs_fraction__3[8], xbs_fraction__3[9], xbs_fraction__3[10], xbs_fraction__3[11], xbs_fraction__3[12], xbs_fraction__3[13], xbs_fraction__3[14], xbs_fraction__3[15], xbs_fraction__3[16], xbs_fraction__3[17], xbs_fraction__3[18], xbs_fraction__3[19], xbs_fraction__3[20], xbs_fraction__3[21], xbs_fraction__3[22], xbs_fraction__3[23], xbs_fraction__3[24], xbs_fraction__3[25], xbs_fraction__3[26], xbs_fraction__3[27]};
  assign one_hot_161097 = {reverse_161089[27:0] == 28'h000_0000, reverse_161089[27] && reverse_161089[26:0] == 27'h000_0000, reverse_161089[26] && reverse_161089[25:0] == 26'h000_0000, reverse_161089[25] && reverse_161089[24:0] == 25'h000_0000, reverse_161089[24] && reverse_161089[23:0] == 24'h00_0000, reverse_161089[23] && reverse_161089[22:0] == 23'h00_0000, reverse_161089[22] && reverse_161089[21:0] == 22'h00_0000, reverse_161089[21] && reverse_161089[20:0] == 21'h00_0000, reverse_161089[20] && reverse_161089[19:0] == 20'h0_0000, reverse_161089[19] && reverse_161089[18:0] == 19'h0_0000, reverse_161089[18] && reverse_161089[17:0] == 18'h0_0000, reverse_161089[17] && reverse_161089[16:0] == 17'h0_0000, reverse_161089[16] && reverse_161089[15:0] == 16'h0000, reverse_161089[15] && reverse_161089[14:0] == 15'h0000, reverse_161089[14] && reverse_161089[13:0] == 14'h0000, reverse_161089[13] && reverse_161089[12:0] == 13'h0000, reverse_161089[12] && reverse_161089[11:0] == 12'h000, reverse_161089[11] && reverse_161089[10:0] == 11'h000, reverse_161089[10] && reverse_161089[9:0] == 10'h000, reverse_161089[9] && reverse_161089[8:0] == 9'h000, reverse_161089[8] && reverse_161089[7:0] == 8'h00, reverse_161089[7] && reverse_161089[6:0] == 7'h00, reverse_161089[6] && reverse_161089[5:0] == 6'h00, reverse_161089[5] && reverse_161089[4:0] == 5'h00, reverse_161089[4] && reverse_161089[3:0] == 4'h0, reverse_161089[3] && reverse_161089[2:0] == 3'h0, reverse_161089[2] && reverse_161089[1:0] == 2'h0, reverse_161089[1] && !reverse_161089[0], reverse_161089[0]};
  assign reverse_161098 = {xbs_fraction__24[0], xbs_fraction__24[1], xbs_fraction__24[2], xbs_fraction__24[3], xbs_fraction__24[4], xbs_fraction__24[5], xbs_fraction__24[6], xbs_fraction__24[7], xbs_fraction__24[8], xbs_fraction__24[9], xbs_fraction__24[10], xbs_fraction__24[11], xbs_fraction__24[12], xbs_fraction__24[13], xbs_fraction__24[14], xbs_fraction__24[15], xbs_fraction__24[16], xbs_fraction__24[17], xbs_fraction__24[18], xbs_fraction__24[19], xbs_fraction__24[20], xbs_fraction__24[21], xbs_fraction__24[22], xbs_fraction__24[23], xbs_fraction__24[24], xbs_fraction__24[25], xbs_fraction__24[26], xbs_fraction__24[27]};
  assign one_hot_161099 = {reverse_161091[27:0] == 28'h000_0000, reverse_161091[27] && reverse_161091[26:0] == 27'h000_0000, reverse_161091[26] && reverse_161091[25:0] == 26'h000_0000, reverse_161091[25] && reverse_161091[24:0] == 25'h000_0000, reverse_161091[24] && reverse_161091[23:0] == 24'h00_0000, reverse_161091[23] && reverse_161091[22:0] == 23'h00_0000, reverse_161091[22] && reverse_161091[21:0] == 22'h00_0000, reverse_161091[21] && reverse_161091[20:0] == 21'h00_0000, reverse_161091[20] && reverse_161091[19:0] == 20'h0_0000, reverse_161091[19] && reverse_161091[18:0] == 19'h0_0000, reverse_161091[18] && reverse_161091[17:0] == 18'h0_0000, reverse_161091[17] && reverse_161091[16:0] == 17'h0_0000, reverse_161091[16] && reverse_161091[15:0] == 16'h0000, reverse_161091[15] && reverse_161091[14:0] == 15'h0000, reverse_161091[14] && reverse_161091[13:0] == 14'h0000, reverse_161091[13] && reverse_161091[12:0] == 13'h0000, reverse_161091[12] && reverse_161091[11:0] == 12'h000, reverse_161091[11] && reverse_161091[10:0] == 11'h000, reverse_161091[10] && reverse_161091[9:0] == 10'h000, reverse_161091[9] && reverse_161091[8:0] == 9'h000, reverse_161091[8] && reverse_161091[7:0] == 8'h00, reverse_161091[7] && reverse_161091[6:0] == 7'h00, reverse_161091[6] && reverse_161091[5:0] == 6'h00, reverse_161091[5] && reverse_161091[4:0] == 5'h00, reverse_161091[4] && reverse_161091[3:0] == 4'h0, reverse_161091[3] && reverse_161091[2:0] == 3'h0, reverse_161091[2] && reverse_161091[1:0] == 2'h0, reverse_161091[1] && !reverse_161091[0], reverse_161091[0]};
  assign reverse_161100 = {xbs_fraction__42[0], xbs_fraction__42[1], xbs_fraction__42[2], xbs_fraction__42[3], xbs_fraction__42[4], xbs_fraction__42[5], xbs_fraction__42[6], xbs_fraction__42[7], xbs_fraction__42[8], xbs_fraction__42[9], xbs_fraction__42[10], xbs_fraction__42[11], xbs_fraction__42[12], xbs_fraction__42[13], xbs_fraction__42[14], xbs_fraction__42[15], xbs_fraction__42[16], xbs_fraction__42[17], xbs_fraction__42[18], xbs_fraction__42[19], xbs_fraction__42[20], xbs_fraction__42[21], xbs_fraction__42[22], xbs_fraction__42[23], xbs_fraction__42[24], xbs_fraction__42[25], xbs_fraction__42[26], xbs_fraction__42[27]};
  assign one_hot_161101 = {reverse_161093[27:0] == 28'h000_0000, reverse_161093[27] && reverse_161093[26:0] == 27'h000_0000, reverse_161093[26] && reverse_161093[25:0] == 26'h000_0000, reverse_161093[25] && reverse_161093[24:0] == 25'h000_0000, reverse_161093[24] && reverse_161093[23:0] == 24'h00_0000, reverse_161093[23] && reverse_161093[22:0] == 23'h00_0000, reverse_161093[22] && reverse_161093[21:0] == 22'h00_0000, reverse_161093[21] && reverse_161093[20:0] == 21'h00_0000, reverse_161093[20] && reverse_161093[19:0] == 20'h0_0000, reverse_161093[19] && reverse_161093[18:0] == 19'h0_0000, reverse_161093[18] && reverse_161093[17:0] == 18'h0_0000, reverse_161093[17] && reverse_161093[16:0] == 17'h0_0000, reverse_161093[16] && reverse_161093[15:0] == 16'h0000, reverse_161093[15] && reverse_161093[14:0] == 15'h0000, reverse_161093[14] && reverse_161093[13:0] == 14'h0000, reverse_161093[13] && reverse_161093[12:0] == 13'h0000, reverse_161093[12] && reverse_161093[11:0] == 12'h000, reverse_161093[11] && reverse_161093[10:0] == 11'h000, reverse_161093[10] && reverse_161093[9:0] == 10'h000, reverse_161093[9] && reverse_161093[8:0] == 9'h000, reverse_161093[8] && reverse_161093[7:0] == 8'h00, reverse_161093[7] && reverse_161093[6:0] == 7'h00, reverse_161093[6] && reverse_161093[5:0] == 6'h00, reverse_161093[5] && reverse_161093[4:0] == 5'h00, reverse_161093[4] && reverse_161093[3:0] == 4'h0, reverse_161093[3] && reverse_161093[2:0] == 3'h0, reverse_161093[2] && reverse_161093[1:0] == 2'h0, reverse_161093[1] && !reverse_161093[0], reverse_161093[0]};
  assign reverse_161102 = {xbs_fraction__60[0], xbs_fraction__60[1], xbs_fraction__60[2], xbs_fraction__60[3], xbs_fraction__60[4], xbs_fraction__60[5], xbs_fraction__60[6], xbs_fraction__60[7], xbs_fraction__60[8], xbs_fraction__60[9], xbs_fraction__60[10], xbs_fraction__60[11], xbs_fraction__60[12], xbs_fraction__60[13], xbs_fraction__60[14], xbs_fraction__60[15], xbs_fraction__60[16], xbs_fraction__60[17], xbs_fraction__60[18], xbs_fraction__60[19], xbs_fraction__60[20], xbs_fraction__60[21], xbs_fraction__60[22], xbs_fraction__60[23], xbs_fraction__60[24], xbs_fraction__60[25], xbs_fraction__60[26], xbs_fraction__60[27]};
  assign one_hot_161103 = {reverse_161095[27:0] == 28'h000_0000, reverse_161095[27] && reverse_161095[26:0] == 27'h000_0000, reverse_161095[26] && reverse_161095[25:0] == 26'h000_0000, reverse_161095[25] && reverse_161095[24:0] == 25'h000_0000, reverse_161095[24] && reverse_161095[23:0] == 24'h00_0000, reverse_161095[23] && reverse_161095[22:0] == 23'h00_0000, reverse_161095[22] && reverse_161095[21:0] == 22'h00_0000, reverse_161095[21] && reverse_161095[20:0] == 21'h00_0000, reverse_161095[20] && reverse_161095[19:0] == 20'h0_0000, reverse_161095[19] && reverse_161095[18:0] == 19'h0_0000, reverse_161095[18] && reverse_161095[17:0] == 18'h0_0000, reverse_161095[17] && reverse_161095[16:0] == 17'h0_0000, reverse_161095[16] && reverse_161095[15:0] == 16'h0000, reverse_161095[15] && reverse_161095[14:0] == 15'h0000, reverse_161095[14] && reverse_161095[13:0] == 14'h0000, reverse_161095[13] && reverse_161095[12:0] == 13'h0000, reverse_161095[12] && reverse_161095[11:0] == 12'h000, reverse_161095[11] && reverse_161095[10:0] == 11'h000, reverse_161095[10] && reverse_161095[9:0] == 10'h000, reverse_161095[9] && reverse_161095[8:0] == 9'h000, reverse_161095[8] && reverse_161095[7:0] == 8'h00, reverse_161095[7] && reverse_161095[6:0] == 7'h00, reverse_161095[6] && reverse_161095[5:0] == 6'h00, reverse_161095[5] && reverse_161095[4:0] == 5'h00, reverse_161095[4] && reverse_161095[3:0] == 4'h0, reverse_161095[3] && reverse_161095[2:0] == 3'h0, reverse_161095[2] && reverse_161095[1:0] == 2'h0, reverse_161095[1] && !reverse_161095[0], reverse_161095[0]};
  assign one_hot_161104 = {reverse_161096[27:0] == 28'h000_0000, reverse_161096[27] && reverse_161096[26:0] == 27'h000_0000, reverse_161096[26] && reverse_161096[25:0] == 26'h000_0000, reverse_161096[25] && reverse_161096[24:0] == 25'h000_0000, reverse_161096[24] && reverse_161096[23:0] == 24'h00_0000, reverse_161096[23] && reverse_161096[22:0] == 23'h00_0000, reverse_161096[22] && reverse_161096[21:0] == 22'h00_0000, reverse_161096[21] && reverse_161096[20:0] == 21'h00_0000, reverse_161096[20] && reverse_161096[19:0] == 20'h0_0000, reverse_161096[19] && reverse_161096[18:0] == 19'h0_0000, reverse_161096[18] && reverse_161096[17:0] == 18'h0_0000, reverse_161096[17] && reverse_161096[16:0] == 17'h0_0000, reverse_161096[16] && reverse_161096[15:0] == 16'h0000, reverse_161096[15] && reverse_161096[14:0] == 15'h0000, reverse_161096[14] && reverse_161096[13:0] == 14'h0000, reverse_161096[13] && reverse_161096[12:0] == 13'h0000, reverse_161096[12] && reverse_161096[11:0] == 12'h000, reverse_161096[11] && reverse_161096[10:0] == 11'h000, reverse_161096[10] && reverse_161096[9:0] == 10'h000, reverse_161096[9] && reverse_161096[8:0] == 9'h000, reverse_161096[8] && reverse_161096[7:0] == 8'h00, reverse_161096[7] && reverse_161096[6:0] == 7'h00, reverse_161096[6] && reverse_161096[5:0] == 6'h00, reverse_161096[5] && reverse_161096[4:0] == 5'h00, reverse_161096[4] && reverse_161096[3:0] == 4'h0, reverse_161096[3] && reverse_161096[2:0] == 3'h0, reverse_161096[2] && reverse_161096[1:0] == 2'h0, reverse_161096[1] && !reverse_161096[0], reverse_161096[0]};
  assign encode_161105 = {one_hot_161097[16] | one_hot_161097[17] | one_hot_161097[18] | one_hot_161097[19] | one_hot_161097[20] | one_hot_161097[21] | one_hot_161097[22] | one_hot_161097[23] | one_hot_161097[24] | one_hot_161097[25] | one_hot_161097[26] | one_hot_161097[27] | one_hot_161097[28], one_hot_161097[8] | one_hot_161097[9] | one_hot_161097[10] | one_hot_161097[11] | one_hot_161097[12] | one_hot_161097[13] | one_hot_161097[14] | one_hot_161097[15] | one_hot_161097[24] | one_hot_161097[25] | one_hot_161097[26] | one_hot_161097[27] | one_hot_161097[28], one_hot_161097[4] | one_hot_161097[5] | one_hot_161097[6] | one_hot_161097[7] | one_hot_161097[12] | one_hot_161097[13] | one_hot_161097[14] | one_hot_161097[15] | one_hot_161097[20] | one_hot_161097[21] | one_hot_161097[22] | one_hot_161097[23] | one_hot_161097[28], one_hot_161097[2] | one_hot_161097[3] | one_hot_161097[6] | one_hot_161097[7] | one_hot_161097[10] | one_hot_161097[11] | one_hot_161097[14] | one_hot_161097[15] | one_hot_161097[18] | one_hot_161097[19] | one_hot_161097[22] | one_hot_161097[23] | one_hot_161097[26] | one_hot_161097[27], one_hot_161097[1] | one_hot_161097[3] | one_hot_161097[5] | one_hot_161097[7] | one_hot_161097[9] | one_hot_161097[11] | one_hot_161097[13] | one_hot_161097[15] | one_hot_161097[17] | one_hot_161097[19] | one_hot_161097[21] | one_hot_161097[23] | one_hot_161097[25] | one_hot_161097[27]};
  assign one_hot_161106 = {reverse_161098[27:0] == 28'h000_0000, reverse_161098[27] && reverse_161098[26:0] == 27'h000_0000, reverse_161098[26] && reverse_161098[25:0] == 26'h000_0000, reverse_161098[25] && reverse_161098[24:0] == 25'h000_0000, reverse_161098[24] && reverse_161098[23:0] == 24'h00_0000, reverse_161098[23] && reverse_161098[22:0] == 23'h00_0000, reverse_161098[22] && reverse_161098[21:0] == 22'h00_0000, reverse_161098[21] && reverse_161098[20:0] == 21'h00_0000, reverse_161098[20] && reverse_161098[19:0] == 20'h0_0000, reverse_161098[19] && reverse_161098[18:0] == 19'h0_0000, reverse_161098[18] && reverse_161098[17:0] == 18'h0_0000, reverse_161098[17] && reverse_161098[16:0] == 17'h0_0000, reverse_161098[16] && reverse_161098[15:0] == 16'h0000, reverse_161098[15] && reverse_161098[14:0] == 15'h0000, reverse_161098[14] && reverse_161098[13:0] == 14'h0000, reverse_161098[13] && reverse_161098[12:0] == 13'h0000, reverse_161098[12] && reverse_161098[11:0] == 12'h000, reverse_161098[11] && reverse_161098[10:0] == 11'h000, reverse_161098[10] && reverse_161098[9:0] == 10'h000, reverse_161098[9] && reverse_161098[8:0] == 9'h000, reverse_161098[8] && reverse_161098[7:0] == 8'h00, reverse_161098[7] && reverse_161098[6:0] == 7'h00, reverse_161098[6] && reverse_161098[5:0] == 6'h00, reverse_161098[5] && reverse_161098[4:0] == 5'h00, reverse_161098[4] && reverse_161098[3:0] == 4'h0, reverse_161098[3] && reverse_161098[2:0] == 3'h0, reverse_161098[2] && reverse_161098[1:0] == 2'h0, reverse_161098[1] && !reverse_161098[0], reverse_161098[0]};
  assign encode_161107 = {one_hot_161099[16] | one_hot_161099[17] | one_hot_161099[18] | one_hot_161099[19] | one_hot_161099[20] | one_hot_161099[21] | one_hot_161099[22] | one_hot_161099[23] | one_hot_161099[24] | one_hot_161099[25] | one_hot_161099[26] | one_hot_161099[27] | one_hot_161099[28], one_hot_161099[8] | one_hot_161099[9] | one_hot_161099[10] | one_hot_161099[11] | one_hot_161099[12] | one_hot_161099[13] | one_hot_161099[14] | one_hot_161099[15] | one_hot_161099[24] | one_hot_161099[25] | one_hot_161099[26] | one_hot_161099[27] | one_hot_161099[28], one_hot_161099[4] | one_hot_161099[5] | one_hot_161099[6] | one_hot_161099[7] | one_hot_161099[12] | one_hot_161099[13] | one_hot_161099[14] | one_hot_161099[15] | one_hot_161099[20] | one_hot_161099[21] | one_hot_161099[22] | one_hot_161099[23] | one_hot_161099[28], one_hot_161099[2] | one_hot_161099[3] | one_hot_161099[6] | one_hot_161099[7] | one_hot_161099[10] | one_hot_161099[11] | one_hot_161099[14] | one_hot_161099[15] | one_hot_161099[18] | one_hot_161099[19] | one_hot_161099[22] | one_hot_161099[23] | one_hot_161099[26] | one_hot_161099[27], one_hot_161099[1] | one_hot_161099[3] | one_hot_161099[5] | one_hot_161099[7] | one_hot_161099[9] | one_hot_161099[11] | one_hot_161099[13] | one_hot_161099[15] | one_hot_161099[17] | one_hot_161099[19] | one_hot_161099[21] | one_hot_161099[23] | one_hot_161099[25] | one_hot_161099[27]};
  assign one_hot_161108 = {reverse_161100[27:0] == 28'h000_0000, reverse_161100[27] && reverse_161100[26:0] == 27'h000_0000, reverse_161100[26] && reverse_161100[25:0] == 26'h000_0000, reverse_161100[25] && reverse_161100[24:0] == 25'h000_0000, reverse_161100[24] && reverse_161100[23:0] == 24'h00_0000, reverse_161100[23] && reverse_161100[22:0] == 23'h00_0000, reverse_161100[22] && reverse_161100[21:0] == 22'h00_0000, reverse_161100[21] && reverse_161100[20:0] == 21'h00_0000, reverse_161100[20] && reverse_161100[19:0] == 20'h0_0000, reverse_161100[19] && reverse_161100[18:0] == 19'h0_0000, reverse_161100[18] && reverse_161100[17:0] == 18'h0_0000, reverse_161100[17] && reverse_161100[16:0] == 17'h0_0000, reverse_161100[16] && reverse_161100[15:0] == 16'h0000, reverse_161100[15] && reverse_161100[14:0] == 15'h0000, reverse_161100[14] && reverse_161100[13:0] == 14'h0000, reverse_161100[13] && reverse_161100[12:0] == 13'h0000, reverse_161100[12] && reverse_161100[11:0] == 12'h000, reverse_161100[11] && reverse_161100[10:0] == 11'h000, reverse_161100[10] && reverse_161100[9:0] == 10'h000, reverse_161100[9] && reverse_161100[8:0] == 9'h000, reverse_161100[8] && reverse_161100[7:0] == 8'h00, reverse_161100[7] && reverse_161100[6:0] == 7'h00, reverse_161100[6] && reverse_161100[5:0] == 6'h00, reverse_161100[5] && reverse_161100[4:0] == 5'h00, reverse_161100[4] && reverse_161100[3:0] == 4'h0, reverse_161100[3] && reverse_161100[2:0] == 3'h0, reverse_161100[2] && reverse_161100[1:0] == 2'h0, reverse_161100[1] && !reverse_161100[0], reverse_161100[0]};
  assign encode_161109 = {one_hot_161101[16] | one_hot_161101[17] | one_hot_161101[18] | one_hot_161101[19] | one_hot_161101[20] | one_hot_161101[21] | one_hot_161101[22] | one_hot_161101[23] | one_hot_161101[24] | one_hot_161101[25] | one_hot_161101[26] | one_hot_161101[27] | one_hot_161101[28], one_hot_161101[8] | one_hot_161101[9] | one_hot_161101[10] | one_hot_161101[11] | one_hot_161101[12] | one_hot_161101[13] | one_hot_161101[14] | one_hot_161101[15] | one_hot_161101[24] | one_hot_161101[25] | one_hot_161101[26] | one_hot_161101[27] | one_hot_161101[28], one_hot_161101[4] | one_hot_161101[5] | one_hot_161101[6] | one_hot_161101[7] | one_hot_161101[12] | one_hot_161101[13] | one_hot_161101[14] | one_hot_161101[15] | one_hot_161101[20] | one_hot_161101[21] | one_hot_161101[22] | one_hot_161101[23] | one_hot_161101[28], one_hot_161101[2] | one_hot_161101[3] | one_hot_161101[6] | one_hot_161101[7] | one_hot_161101[10] | one_hot_161101[11] | one_hot_161101[14] | one_hot_161101[15] | one_hot_161101[18] | one_hot_161101[19] | one_hot_161101[22] | one_hot_161101[23] | one_hot_161101[26] | one_hot_161101[27], one_hot_161101[1] | one_hot_161101[3] | one_hot_161101[5] | one_hot_161101[7] | one_hot_161101[9] | one_hot_161101[11] | one_hot_161101[13] | one_hot_161101[15] | one_hot_161101[17] | one_hot_161101[19] | one_hot_161101[21] | one_hot_161101[23] | one_hot_161101[25] | one_hot_161101[27]};
  assign one_hot_161110 = {reverse_161102[27:0] == 28'h000_0000, reverse_161102[27] && reverse_161102[26:0] == 27'h000_0000, reverse_161102[26] && reverse_161102[25:0] == 26'h000_0000, reverse_161102[25] && reverse_161102[24:0] == 25'h000_0000, reverse_161102[24] && reverse_161102[23:0] == 24'h00_0000, reverse_161102[23] && reverse_161102[22:0] == 23'h00_0000, reverse_161102[22] && reverse_161102[21:0] == 22'h00_0000, reverse_161102[21] && reverse_161102[20:0] == 21'h00_0000, reverse_161102[20] && reverse_161102[19:0] == 20'h0_0000, reverse_161102[19] && reverse_161102[18:0] == 19'h0_0000, reverse_161102[18] && reverse_161102[17:0] == 18'h0_0000, reverse_161102[17] && reverse_161102[16:0] == 17'h0_0000, reverse_161102[16] && reverse_161102[15:0] == 16'h0000, reverse_161102[15] && reverse_161102[14:0] == 15'h0000, reverse_161102[14] && reverse_161102[13:0] == 14'h0000, reverse_161102[13] && reverse_161102[12:0] == 13'h0000, reverse_161102[12] && reverse_161102[11:0] == 12'h000, reverse_161102[11] && reverse_161102[10:0] == 11'h000, reverse_161102[10] && reverse_161102[9:0] == 10'h000, reverse_161102[9] && reverse_161102[8:0] == 9'h000, reverse_161102[8] && reverse_161102[7:0] == 8'h00, reverse_161102[7] && reverse_161102[6:0] == 7'h00, reverse_161102[6] && reverse_161102[5:0] == 6'h00, reverse_161102[5] && reverse_161102[4:0] == 5'h00, reverse_161102[4] && reverse_161102[3:0] == 4'h0, reverse_161102[3] && reverse_161102[2:0] == 3'h0, reverse_161102[2] && reverse_161102[1:0] == 2'h0, reverse_161102[1] && !reverse_161102[0], reverse_161102[0]};
  assign encode_161111 = {one_hot_161103[16] | one_hot_161103[17] | one_hot_161103[18] | one_hot_161103[19] | one_hot_161103[20] | one_hot_161103[21] | one_hot_161103[22] | one_hot_161103[23] | one_hot_161103[24] | one_hot_161103[25] | one_hot_161103[26] | one_hot_161103[27] | one_hot_161103[28], one_hot_161103[8] | one_hot_161103[9] | one_hot_161103[10] | one_hot_161103[11] | one_hot_161103[12] | one_hot_161103[13] | one_hot_161103[14] | one_hot_161103[15] | one_hot_161103[24] | one_hot_161103[25] | one_hot_161103[26] | one_hot_161103[27] | one_hot_161103[28], one_hot_161103[4] | one_hot_161103[5] | one_hot_161103[6] | one_hot_161103[7] | one_hot_161103[12] | one_hot_161103[13] | one_hot_161103[14] | one_hot_161103[15] | one_hot_161103[20] | one_hot_161103[21] | one_hot_161103[22] | one_hot_161103[23] | one_hot_161103[28], one_hot_161103[2] | one_hot_161103[3] | one_hot_161103[6] | one_hot_161103[7] | one_hot_161103[10] | one_hot_161103[11] | one_hot_161103[14] | one_hot_161103[15] | one_hot_161103[18] | one_hot_161103[19] | one_hot_161103[22] | one_hot_161103[23] | one_hot_161103[26] | one_hot_161103[27], one_hot_161103[1] | one_hot_161103[3] | one_hot_161103[5] | one_hot_161103[7] | one_hot_161103[9] | one_hot_161103[11] | one_hot_161103[13] | one_hot_161103[15] | one_hot_161103[17] | one_hot_161103[19] | one_hot_161103[21] | one_hot_161103[23] | one_hot_161103[25] | one_hot_161103[27]};
  assign encode_161112 = {one_hot_161104[16] | one_hot_161104[17] | one_hot_161104[18] | one_hot_161104[19] | one_hot_161104[20] | one_hot_161104[21] | one_hot_161104[22] | one_hot_161104[23] | one_hot_161104[24] | one_hot_161104[25] | one_hot_161104[26] | one_hot_161104[27] | one_hot_161104[28], one_hot_161104[8] | one_hot_161104[9] | one_hot_161104[10] | one_hot_161104[11] | one_hot_161104[12] | one_hot_161104[13] | one_hot_161104[14] | one_hot_161104[15] | one_hot_161104[24] | one_hot_161104[25] | one_hot_161104[26] | one_hot_161104[27] | one_hot_161104[28], one_hot_161104[4] | one_hot_161104[5] | one_hot_161104[6] | one_hot_161104[7] | one_hot_161104[12] | one_hot_161104[13] | one_hot_161104[14] | one_hot_161104[15] | one_hot_161104[20] | one_hot_161104[21] | one_hot_161104[22] | one_hot_161104[23] | one_hot_161104[28], one_hot_161104[2] | one_hot_161104[3] | one_hot_161104[6] | one_hot_161104[7] | one_hot_161104[10] | one_hot_161104[11] | one_hot_161104[14] | one_hot_161104[15] | one_hot_161104[18] | one_hot_161104[19] | one_hot_161104[22] | one_hot_161104[23] | one_hot_161104[26] | one_hot_161104[27], one_hot_161104[1] | one_hot_161104[3] | one_hot_161104[5] | one_hot_161104[7] | one_hot_161104[9] | one_hot_161104[11] | one_hot_161104[13] | one_hot_161104[15] | one_hot_161104[17] | one_hot_161104[19] | one_hot_161104[21] | one_hot_161104[23] | one_hot_161104[25] | one_hot_161104[27]};
  assign encode_161114 = {one_hot_161106[16] | one_hot_161106[17] | one_hot_161106[18] | one_hot_161106[19] | one_hot_161106[20] | one_hot_161106[21] | one_hot_161106[22] | one_hot_161106[23] | one_hot_161106[24] | one_hot_161106[25] | one_hot_161106[26] | one_hot_161106[27] | one_hot_161106[28], one_hot_161106[8] | one_hot_161106[9] | one_hot_161106[10] | one_hot_161106[11] | one_hot_161106[12] | one_hot_161106[13] | one_hot_161106[14] | one_hot_161106[15] | one_hot_161106[24] | one_hot_161106[25] | one_hot_161106[26] | one_hot_161106[27] | one_hot_161106[28], one_hot_161106[4] | one_hot_161106[5] | one_hot_161106[6] | one_hot_161106[7] | one_hot_161106[12] | one_hot_161106[13] | one_hot_161106[14] | one_hot_161106[15] | one_hot_161106[20] | one_hot_161106[21] | one_hot_161106[22] | one_hot_161106[23] | one_hot_161106[28], one_hot_161106[2] | one_hot_161106[3] | one_hot_161106[6] | one_hot_161106[7] | one_hot_161106[10] | one_hot_161106[11] | one_hot_161106[14] | one_hot_161106[15] | one_hot_161106[18] | one_hot_161106[19] | one_hot_161106[22] | one_hot_161106[23] | one_hot_161106[26] | one_hot_161106[27], one_hot_161106[1] | one_hot_161106[3] | one_hot_161106[5] | one_hot_161106[7] | one_hot_161106[9] | one_hot_161106[11] | one_hot_161106[13] | one_hot_161106[15] | one_hot_161106[17] | one_hot_161106[19] | one_hot_161106[21] | one_hot_161106[23] | one_hot_161106[25] | one_hot_161106[27]};
  assign encode_161116 = {one_hot_161108[16] | one_hot_161108[17] | one_hot_161108[18] | one_hot_161108[19] | one_hot_161108[20] | one_hot_161108[21] | one_hot_161108[22] | one_hot_161108[23] | one_hot_161108[24] | one_hot_161108[25] | one_hot_161108[26] | one_hot_161108[27] | one_hot_161108[28], one_hot_161108[8] | one_hot_161108[9] | one_hot_161108[10] | one_hot_161108[11] | one_hot_161108[12] | one_hot_161108[13] | one_hot_161108[14] | one_hot_161108[15] | one_hot_161108[24] | one_hot_161108[25] | one_hot_161108[26] | one_hot_161108[27] | one_hot_161108[28], one_hot_161108[4] | one_hot_161108[5] | one_hot_161108[6] | one_hot_161108[7] | one_hot_161108[12] | one_hot_161108[13] | one_hot_161108[14] | one_hot_161108[15] | one_hot_161108[20] | one_hot_161108[21] | one_hot_161108[22] | one_hot_161108[23] | one_hot_161108[28], one_hot_161108[2] | one_hot_161108[3] | one_hot_161108[6] | one_hot_161108[7] | one_hot_161108[10] | one_hot_161108[11] | one_hot_161108[14] | one_hot_161108[15] | one_hot_161108[18] | one_hot_161108[19] | one_hot_161108[22] | one_hot_161108[23] | one_hot_161108[26] | one_hot_161108[27], one_hot_161108[1] | one_hot_161108[3] | one_hot_161108[5] | one_hot_161108[7] | one_hot_161108[9] | one_hot_161108[11] | one_hot_161108[13] | one_hot_161108[15] | one_hot_161108[17] | one_hot_161108[19] | one_hot_161108[21] | one_hot_161108[23] | one_hot_161108[25] | one_hot_161108[27]};
  assign encode_161118 = {one_hot_161110[16] | one_hot_161110[17] | one_hot_161110[18] | one_hot_161110[19] | one_hot_161110[20] | one_hot_161110[21] | one_hot_161110[22] | one_hot_161110[23] | one_hot_161110[24] | one_hot_161110[25] | one_hot_161110[26] | one_hot_161110[27] | one_hot_161110[28], one_hot_161110[8] | one_hot_161110[9] | one_hot_161110[10] | one_hot_161110[11] | one_hot_161110[12] | one_hot_161110[13] | one_hot_161110[14] | one_hot_161110[15] | one_hot_161110[24] | one_hot_161110[25] | one_hot_161110[26] | one_hot_161110[27] | one_hot_161110[28], one_hot_161110[4] | one_hot_161110[5] | one_hot_161110[6] | one_hot_161110[7] | one_hot_161110[12] | one_hot_161110[13] | one_hot_161110[14] | one_hot_161110[15] | one_hot_161110[20] | one_hot_161110[21] | one_hot_161110[22] | one_hot_161110[23] | one_hot_161110[28], one_hot_161110[2] | one_hot_161110[3] | one_hot_161110[6] | one_hot_161110[7] | one_hot_161110[10] | one_hot_161110[11] | one_hot_161110[14] | one_hot_161110[15] | one_hot_161110[18] | one_hot_161110[19] | one_hot_161110[22] | one_hot_161110[23] | one_hot_161110[26] | one_hot_161110[27], one_hot_161110[1] | one_hot_161110[3] | one_hot_161110[5] | one_hot_161110[7] | one_hot_161110[9] | one_hot_161110[11] | one_hot_161110[13] | one_hot_161110[15] | one_hot_161110[17] | one_hot_161110[19] | one_hot_161110[21] | one_hot_161110[23] | one_hot_161110[25] | one_hot_161110[27]};
  assign cancel__12 = |encode_161105[4:1];
  assign carry_bit__11 = xbs_fraction__11[27];
  assign result_fraction__490 = 23'h00_0000;
  assign cancel__24 = |encode_161107[4:1];
  assign carry_bit__24 = xbs_fraction__23[27];
  assign result_fraction__557 = 23'h00_0000;
  assign cancel__43 = |encode_161109[4:1];
  assign carry_bit__43 = xbs_fraction__41[27];
  assign result_fraction__620 = 23'h00_0000;
  assign cancel__62 = |encode_161111[4:1];
  assign carry_bit__62 = xbs_fraction__59[27];
  assign result_fraction__691 = 23'h00_0000;
  assign cancel__3 = |encode_161112[4:1];
  assign carry_bit__3 = xbs_fraction__3[27];
  assign result_fraction__491 = 23'h00_0000;
  assign leading_zeroes__11 = {result_fraction__490, encode_161105};
  assign cancel__25 = |encode_161114[4:1];
  assign carry_bit__25 = xbs_fraction__24[27];
  assign result_fraction__558 = 23'h00_0000;
  assign leading_zeroes__24 = {result_fraction__557, encode_161107};
  assign cancel__44 = |encode_161116[4:1];
  assign carry_bit__44 = xbs_fraction__42[27];
  assign result_fraction__621 = 23'h00_0000;
  assign leading_zeroes__43 = {result_fraction__620, encode_161109};
  assign cancel__63 = |encode_161118[4:1];
  assign carry_bit__63 = xbs_fraction__60[27];
  assign result_fraction__692 = 23'h00_0000;
  assign leading_zeroes__62 = {result_fraction__691, encode_161111};
  assign leading_zeroes__3 = {result_fraction__491, encode_161112};
  assign carry_fraction__22 = xbs_fraction__11[27:1];
  assign add_161186 = leading_zeroes__11 + 28'hfff_ffff;
  assign leading_zeroes__25 = {result_fraction__558, encode_161114};
  assign carry_fraction__47 = xbs_fraction__23[27:1];
  assign add_161199 = leading_zeroes__24 + 28'hfff_ffff;
  assign leading_zeroes__44 = {result_fraction__621, encode_161116};
  assign array_index_161206 = in_img_unflattened[4'h8];
  assign carry_fraction__85 = xbs_fraction__41[27:1];
  assign add_161213 = leading_zeroes__43 + 28'hfff_ffff;
  assign leading_zeroes__63 = {result_fraction__692, encode_161118};
  assign array_index_161220 = in_img_unflattened[4'h9];
  assign carry_fraction__123 = xbs_fraction__59[27:1];
  assign add_161227 = leading_zeroes__62 + 28'hfff_ffff;
  assign carry_fraction__5 = xbs_fraction__3[27:1];
  assign add_161234 = leading_zeroes__3 + 28'hfff_ffff;
  assign concat_161235 = {~(carry_bit__11 | cancel__12), ~(carry_bit__11 | ~cancel__12), ~(~carry_bit__11 | cancel__12)};
  assign carry_fraction__23 = carry_fraction__22 | {26'h000_0000, xbs_fraction__11[0]};
  assign cancel_fraction__11 = add_161186 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__11[26:0] << add_161186;
  assign carry_fraction__48 = xbs_fraction__24[27:1];
  assign add_161244 = leading_zeroes__25 + 28'hfff_ffff;
  assign concat_161245 = {~(carry_bit__24 | cancel__24), ~(carry_bit__24 | ~cancel__24), ~(~carry_bit__24 | cancel__24)};
  assign carry_fraction__49 = carry_fraction__47 | {26'h000_0000, xbs_fraction__23[0]};
  assign cancel_fraction__24 = add_161199 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__23[26:0] << add_161199;
  assign carry_fraction__86 = xbs_fraction__42[27:1];
  assign add_161254 = leading_zeroes__44 + 28'hfff_ffff;
  assign x_bexp__334 = array_index_161206[30:23];
  assign concat_161256 = {~(carry_bit__43 | cancel__43), ~(carry_bit__43 | ~cancel__43), ~(~carry_bit__43 | cancel__43)};
  assign carry_fraction__87 = carry_fraction__85 | {26'h000_0000, xbs_fraction__41[0]};
  assign cancel_fraction__43 = add_161213 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__41[26:0] << add_161213;
  assign carry_fraction__124 = xbs_fraction__60[27:1];
  assign add_161265 = leading_zeroes__63 + 28'hfff_ffff;
  assign x_bexp__478 = array_index_161220[30:23];
  assign concat_161267 = {~(carry_bit__62 | cancel__62), ~(carry_bit__62 | ~cancel__62), ~(~carry_bit__62 | cancel__62)};
  assign carry_fraction__125 = carry_fraction__123 | {26'h000_0000, xbs_fraction__59[0]};
  assign cancel_fraction__62 = add_161227 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__59[26:0] << add_161227;
  assign concat_161270 = {~(carry_bit__3 | cancel__3), ~(carry_bit__3 | ~cancel__3), ~(~carry_bit__3 | cancel__3)};
  assign carry_fraction__6 = carry_fraction__5 | {26'h000_0000, xbs_fraction__3[0]};
  assign cancel_fraction__3 = add_161234 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__3[26:0] << add_161234;
  assign result_sign__988 = 1'h0;
  assign shifted_fraction__11 = carry_fraction__23 & {27{concat_161235[0]}} | cancel_fraction__11 & {27{concat_161235[1]}} | xbs_fraction__11[26:0] & {27{concat_161235[2]}};
  assign concat_161276 = {~(carry_bit__25 | cancel__25), ~(carry_bit__25 | ~cancel__25), ~(~carry_bit__25 | cancel__25)};
  assign carry_fraction__50 = carry_fraction__48 | {26'h000_0000, xbs_fraction__24[0]};
  assign cancel_fraction__25 = add_161244 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__24[26:0] << add_161244;
  assign shifted_fraction__24 = carry_fraction__49 & {27{concat_161245[0]}} | cancel_fraction__24 & {27{concat_161245[1]}} | xbs_fraction__23[26:0] & {27{concat_161245[2]}};
  assign concat_161280 = {~(carry_bit__44 | cancel__44), ~(carry_bit__44 | ~cancel__44), ~(~carry_bit__44 | cancel__44)};
  assign carry_fraction__88 = carry_fraction__86 | {26'h000_0000, xbs_fraction__42[0]};
  assign cancel_fraction__44 = add_161254 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__42[26:0] << add_161254;
  assign result_sign__989 = 1'h0;
  assign shifted_fraction__43 = carry_fraction__87 & {27{concat_161256[0]}} | cancel_fraction__43 & {27{concat_161256[1]}} | xbs_fraction__41[26:0] & {27{concat_161256[2]}};
  assign concat_161286 = {~(carry_bit__63 | cancel__63), ~(carry_bit__63 | ~cancel__63), ~(~carry_bit__63 | cancel__63)};
  assign carry_fraction__126 = carry_fraction__124 | {26'h000_0000, xbs_fraction__60[0]};
  assign cancel_fraction__63 = add_161265 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__60[26:0] << add_161265;
  assign result_sign__990 = 1'h0;
  assign shifted_fraction__62 = carry_fraction__125 & {27{concat_161267[0]}} | cancel_fraction__62 & {27{concat_161267[1]}} | xbs_fraction__59[26:0] & {27{concat_161267[2]}};
  assign shifted_fraction__3 = carry_fraction__6 & {27{concat_161270[0]}} | cancel_fraction__3 & {27{concat_161270[1]}} | xbs_fraction__3[26:0] & {27{concat_161270[2]}};
  assign result_sign__991 = 1'h0;
  assign shifted_fraction__25 = carry_fraction__50 & {27{concat_161276[0]}} | cancel_fraction__25 & {27{concat_161276[1]}} | xbs_fraction__24[26:0] & {27{concat_161276[2]}};
  assign result_sign__992 = 1'h0;
  assign shifted_fraction__44 = carry_fraction__88 & {27{concat_161280[0]}} | cancel_fraction__44 & {27{concat_161280[1]}} | xbs_fraction__42[26:0] & {27{concat_161280[2]}};
  assign result_sign__993 = 1'h0;
  assign shifted_fraction__63 = carry_fraction__126 & {27{concat_161286[0]}} | cancel_fraction__63 & {27{concat_161286[1]}} | xbs_fraction__60[26:0] & {27{concat_161286[2]}};
  assign result_sign__994 = 1'h0;
  assign result_sign__995 = 1'h0;
  assign result_sign__1105 = 1'h0;
  assign add_161313 = {result_sign__988, x_bexp__289[7]} + 2'h1;
  assign normal_chunk__11 = shifted_fraction__11[2:0];
  assign fraction_shift__233 = 3'h4;
  assign half_way_chunk__11 = shifted_fraction__11[3:2];
  assign result_sign__996 = 1'h0;
  assign normal_chunk__24 = shifted_fraction__24[2:0];
  assign fraction_shift__268 = 3'h4;
  assign half_way_chunk__24 = shifted_fraction__24[3:2];
  assign result_sign__997 = 1'h0;
  assign result_sign__1109 = 1'h0;
  assign add_161332 = {result_sign__989, x_bexp__334[7]} + 2'h1;
  assign x_bexp__708 = 8'h00;
  assign result_sign__598 = 1'h0;
  assign x_fraction__334 = array_index_161206[22:0];
  assign normal_chunk__43 = shifted_fraction__43[2:0];
  assign fraction_shift__303 = 3'h4;
  assign half_way_chunk__43 = shifted_fraction__43[3:2];
  assign result_sign__998 = 1'h0;
  assign result_sign__1113 = 1'h0;
  assign add_161346 = {result_sign__990, x_bexp__478[7]} + 2'h1;
  assign x_bexp__709 = 8'h00;
  assign result_sign__704 = 1'h0;
  assign x_fraction__478 = array_index_161220[22:0];
  assign normal_chunk__62 = shifted_fraction__62[2:0];
  assign fraction_shift__338 = 3'h4;
  assign half_way_chunk__62 = shifted_fraction__62[3:2];
  assign normal_chunk__3 = shifted_fraction__3[2:0];
  assign fraction_shift__234 = 3'h4;
  assign half_way_chunk__3 = shifted_fraction__3[3:2];
  assign result_sign__406 = 1'h0;
  assign add_161368 = {result_sign__991, shifted_fraction__11[26:3]} + 25'h000_0001;
  assign normal_chunk__25 = shifted_fraction__25[2:0];
  assign fraction_shift__269 = 3'h4;
  assign half_way_chunk__25 = shifted_fraction__25[3:2];
  assign result_sign__503 = 1'h0;
  assign add_161378 = {result_sign__992, shifted_fraction__24[26:3]} + 25'h000_0001;
  assign normal_chunk__44 = shifted_fraction__44[2:0];
  assign fraction_shift__304 = 3'h4;
  assign half_way_chunk__44 = shifted_fraction__44[3:2];
  assign ne_161387 = x_bexp__334 != x_bexp__708;
  assign result_sign__596 = 1'h0;
  assign add_161393 = {result_sign__993, shifted_fraction__43[26:3]} + 25'h000_0001;
  assign normal_chunk__63 = shifted_fraction__63[2:0];
  assign fraction_shift__339 = 3'h4;
  assign half_way_chunk__63 = shifted_fraction__63[3:2];
  assign ne_161402 = x_bexp__478 != x_bexp__709;
  assign result_sign__702 = 1'h0;
  assign add_161408 = {result_sign__994, shifted_fraction__62[26:3]} + 25'h000_0001;
  assign result_sign__407 = 1'h0;
  assign add_161412 = {result_sign__995, shifted_fraction__3[26:3]} + 25'h000_0001;
  assign exp__13 = {result_sign__1105, add_161313, x_bexp__289[6:0]} + 10'h381;
  assign do_round_up__23 = normal_chunk__11 > fraction_shift__233 | half_way_chunk__11 == 2'h3;
  assign result_sign__504 = 1'h0;
  assign add_161420 = {result_sign__996, shifted_fraction__25[26:3]} + 25'h000_0001;
  assign do_round_up__50 = normal_chunk__24 > fraction_shift__268 | half_way_chunk__24 == 2'h3;
  assign result_sign__597 = 1'h0;
  assign add_161427 = {result_sign__997, shifted_fraction__44[26:3]} + 25'h000_0001;
  assign exp__190 = {result_sign__1109, add_161332, x_bexp__334[6:0]} + 10'h381;
  assign sign_ext_161429 = {10{ne_161387}};
  assign x_fraction__336 = {result_sign__598, x_fraction__334} | 24'h80_0000;
  assign do_round_up__89 = normal_chunk__43 > fraction_shift__303 | half_way_chunk__43 == 2'h3;
  assign result_sign__703 = 1'h0;
  assign add_161438 = {result_sign__998, shifted_fraction__63[26:3]} + 25'h000_0001;
  assign exp__272 = {result_sign__1113, add_161346, x_bexp__478[6:0]} + 10'h381;
  assign sign_ext_161440 = {10{ne_161402}};
  assign x_fraction__480 = {result_sign__704, x_fraction__478} | 24'h80_0000;
  assign do_round_up__128 = normal_chunk__62 > fraction_shift__338 | half_way_chunk__62 == 2'h3;
  assign do_round_up__6 = normal_chunk__3 > fraction_shift__234 | half_way_chunk__3 == 2'h3;
  assign exp__14 = exp__13 & sign_ext_157981;
  assign rounded_fraction__11 = do_round_up__23 ? {add_161368, normal_chunk__11} : {result_sign__406, shifted_fraction__11};
  assign do_round_up__51 = normal_chunk__25 > fraction_shift__269 | half_way_chunk__25 == 2'h3;
  assign rounded_fraction__24 = do_round_up__50 ? {add_161378, normal_chunk__24} : {result_sign__503, shifted_fraction__24};
  assign do_round_up__90 = normal_chunk__44 > fraction_shift__304 | half_way_chunk__44 == 2'h3;
  assign exp__192 = exp__190 & sign_ext_161429;
  assign x_fraction__338 = x_fraction__336 & {24{ne_161387}};
  assign result_sign__812 = 1'h0;
  assign result_sign__813 = 1'h0;
  assign rounded_fraction__43 = do_round_up__89 ? {add_161393, normal_chunk__43} : {result_sign__596, shifted_fraction__43};
  assign do_round_up__129 = normal_chunk__63 > fraction_shift__339 | half_way_chunk__63 == 2'h3;
  assign exp__274 = exp__272 & sign_ext_161440;
  assign x_fraction__482 = x_fraction__480 & {24{ne_161402}};
  assign result_sign__814 = 1'h0;
  assign result_sign__815 = 1'h0;
  assign rounded_fraction__62 = do_round_up__128 ? {add_161408, normal_chunk__62} : {result_sign__702, shifted_fraction__62};
  assign rounded_fraction__3 = do_round_up__6 ? {add_161412, normal_chunk__3} : {result_sign__407, shifted_fraction__3};
  assign result_sign__408 = 1'h0;
  assign x_bexp__578 = 8'h00;
  assign rounding_carry__11 = rounded_fraction__11[27];
  assign rounded_fraction__25 = do_round_up__51 ? {add_161420, normal_chunk__25} : {result_sign__504, shifted_fraction__25};
  assign result_sign__505 = 1'h0;
  assign x_bexp__596 = 8'h00;
  assign rounding_carry__24 = rounded_fraction__24[27];
  assign rounded_fraction__44 = do_round_up__90 ? {add_161427, normal_chunk__44} : {result_sign__597, shifted_fraction__44};
  assign concat_161485 = {x_fraction__338, result_sign__812};
  assign concat_161486 = {result_sign__813, x_fraction__338};
  assign result_sign__600 = 1'h0;
  assign x_bexp__614 = 8'h00;
  assign rounding_carry__43 = rounded_fraction__43[27];
  assign rounded_fraction__63 = do_round_up__129 ? {add_161438, normal_chunk__63} : {result_sign__703, shifted_fraction__63};
  assign concat_161492 = {x_fraction__482, result_sign__814};
  assign concat_161493 = {result_sign__815, x_fraction__482};
  assign result_sign__706 = 1'h0;
  assign x_bexp__632 = 8'h00;
  assign rounding_carry__62 = rounded_fraction__62[27];
  assign result_sign__409 = 1'h0;
  assign x_bexp__579 = 8'h00;
  assign rounding_carry__3 = rounded_fraction__3[27];
  assign sel_161500 = $signed(exp__14) <= $signed(10'h000) ? concat_158016 : concat_158015;
  assign result_sign__506 = 1'h0;
  assign x_bexp__597 = 8'h00;
  assign rounding_carry__25 = rounded_fraction__25[27];
  assign result_sign__601 = 1'h0;
  assign x_bexp__615 = 8'h00;
  assign rounding_carry__44 = rounded_fraction__44[27];
  assign sel_161511 = $signed(exp__192) <= $signed(10'h000) ? concat_161486 : concat_161485;
  assign result_sign__707 = 1'h0;
  assign x_bexp__633 = 8'h00;
  assign rounding_carry__63 = rounded_fraction__63[27];
  assign sel_161517 = $signed(exp__274) <= $signed(10'h000) ? concat_161493 : concat_161492;
  assign result_sign__931 = 1'h0;
  assign fraction__33 = sel_161500[23:1];
  assign result_sign__410 = 1'h0;
  assign add_161525 = {result_sign__408, x_bexp__94} + {x_bexp__578, rounding_carry__11};
  assign result_sign__507 = 1'h0;
  assign add_161531 = {result_sign__505, x_bexp__187} + {x_bexp__596, rounding_carry__24};
  assign result_sign__943 = 1'h0;
  assign fraction__424 = sel_161511[23:1];
  assign result_sign__602 = 1'h0;
  assign add_161539 = {result_sign__600, x_bexp__331} + {x_bexp__614, rounding_carry__43};
  assign result_sign__951 = 1'h0;
  assign fraction__603 = sel_161517[23:1];
  assign result_sign__708 = 1'h0;
  assign add_161547 = {result_sign__706, x_bexp__475} + {x_bexp__632, rounding_carry__62};
  assign result_sign__411 = 1'h0;
  assign add_161551 = {result_sign__409, x_bexp__22} + {x_bexp__579, rounding_carry__3};
  assign fraction__34 = {result_sign__931, fraction__33};
  assign result_sign__508 = 1'h0;
  assign add_161564 = {result_sign__506, x_bexp__188} + {x_bexp__597, rounding_carry__25};
  assign result_sign__603 = 1'h0;
  assign add_161573 = {result_sign__601, x_bexp__332} + {x_bexp__615, rounding_carry__44};
  assign fraction__426 = {result_sign__943, fraction__424};
  assign result_sign__709 = 1'h0;
  assign add_161586 = {result_sign__707, x_bexp__476} + {x_bexp__633, rounding_carry__63};
  assign fraction__605 = {result_sign__951, fraction__603};
  assign do_round_up__7 = sel_161500[0] & sel_161500[1];
  assign add_161604 = fraction__34 + 24'h00_0001;
  assign add_161605 = {result_sign__410, add_161525} + 10'h001;
  assign add_161613 = {result_sign__507, add_161531} + 10'h001;
  assign do_round_up__92 = sel_161511[0] & sel_161511[1];
  assign add_161622 = fraction__426 + 24'h00_0001;
  assign add_161623 = {result_sign__602, add_161539} + 10'h001;
  assign do_round_up__131 = sel_161517[0] & sel_161517[1];
  assign add_161632 = fraction__605 + 24'h00_0001;
  assign add_161633 = {result_sign__708, add_161547} + 10'h001;
  assign add_161636 = {result_sign__411, add_161551} + 10'h001;
  assign fraction__35 = do_round_up__7 ? add_161604 : fraction__34;
  assign wide_exponent__33 = add_161605 - {5'h00, encode_161105};
  assign add_161643 = {result_sign__508, add_161564} + 10'h001;
  assign wide_exponent__70 = add_161613 - {5'h00, encode_161107};
  assign add_161648 = {result_sign__603, add_161573} + 10'h001;
  assign fraction__428 = do_round_up__92 ? add_161622 : fraction__426;
  assign wide_exponent__127 = add_161623 - {5'h00, encode_161109};
  assign add_161655 = {result_sign__709, add_161586} + 10'h001;
  assign fraction__607 = do_round_up__131 ? add_161632 : fraction__605;
  assign wide_exponent__184 = add_161633 - {5'h00, encode_161111};
  assign wide_exponent__7 = add_161636 - {5'h00, encode_161112};
  assign add_161665 = exp__14 + 10'h001;
  assign wide_exponent__34 = wide_exponent__33 & {10{add_161030 != 26'h000_0000 | xddend_y__11[2:0] != 3'h0}};
  assign wide_exponent__71 = add_161643 - {5'h00, encode_161114};
  assign wide_exponent__72 = wide_exponent__70 & {10{add_161033 != 26'h000_0000 | xddend_y__23[2:0] != 3'h0}};
  assign wide_exponent__128 = add_161648 - {5'h00, encode_161116};
  assign add_161673 = exp__192 + 10'h001;
  assign wide_exponent__129 = wide_exponent__127 & {10{add_161036 != 26'h000_0000 | xddend_y__41[2:0] != 3'h0}};
  assign wide_exponent__185 = add_161655 - {5'h00, encode_161118};
  assign add_161678 = exp__274 + 10'h001;
  assign wide_exponent__186 = wide_exponent__184 & {10{add_161039 != 26'h000_0000 | xddend_y__59[2:0] != 3'h0}};
  assign wide_exponent__8 = wide_exponent__7 & {10{add_161040 != 26'h000_0000 | xddend_y__3[2:0] != 3'h0}};
  assign exp__16 = fraction__35[23] ? add_161665 : exp__14;
  assign high_exp__367 = 8'hff;
  assign result_fraction__773 = 23'h00_0000;
  assign high_exp__368 = 8'hff;
  assign result_fraction__774 = 23'h00_0000;
  assign high_exp__91 = 8'hff;
  assign result_fraction__492 = 23'h00_0000;
  assign high_exp__92 = 8'hff;
  assign result_fraction__493 = 23'h00_0000;
  assign wide_exponent__73 = wide_exponent__71 & {10{add_161043 != 26'h000_0000 | xddend_y__24[2:0] != 3'h0}};
  assign high_exp__399 = 8'hff;
  assign result_fraction__806 = 23'h00_0000;
  assign high_exp__400 = 8'hff;
  assign result_fraction__807 = 23'h00_0000;
  assign high_exp__156 = 8'hff;
  assign result_fraction__559 = 23'h00_0000;
  assign high_exp__157 = 8'hff;
  assign result_fraction__560 = 23'h00_0000;
  assign wide_exponent__130 = wide_exponent__128 & {10{add_161046 != 26'h000_0000 | xddend_y__42[2:0] != 3'h0}};
  assign exp__196 = fraction__428[23] ? add_161673 : exp__192;
  assign high_exp__431 = 8'hff;
  assign result_fraction__839 = 23'h00_0000;
  assign high_exp__432 = 8'hff;
  assign result_fraction__840 = 23'h00_0000;
  assign high_exp__220 = 8'hff;
  assign result_fraction__622 = 23'h00_0000;
  assign high_exp__221 = 8'hff;
  assign result_fraction__623 = 23'h00_0000;
  assign wide_exponent__187 = wide_exponent__185 & {10{add_161049 != 26'h000_0000 | xddend_y__60[2:0] != 3'h0}};
  assign exp__278 = fraction__607[23] ? add_161678 : exp__274;
  assign high_exp__463 = 8'hff;
  assign result_fraction__872 = 23'h00_0000;
  assign high_exp__464 = 8'hff;
  assign result_fraction__873 = 23'h00_0000;
  assign high_exp__290 = 8'hff;
  assign result_fraction__693 = 23'h00_0000;
  assign high_exp__291 = 8'hff;
  assign result_fraction__694 = 23'h00_0000;
  assign high_exp__353 = 8'hff;
  assign result_fraction__758 = 23'h00_0000;
  assign high_exp__354 = 8'hff;
  assign result_fraction__759 = 23'h00_0000;
  assign high_exp__93 = 8'hff;
  assign result_fraction__494 = 23'h00_0000;
  assign high_exp__94 = 8'hff;
  assign result_fraction__495 = 23'h00_0000;
  assign ne_161738 = x_fraction__94 != result_fraction__773;
  assign ne_161740 = prod_fraction__33 != result_fraction__774;
  assign eq_161741 = x_bexp__94 == high_exp__91;
  assign eq_161742 = x_fraction__94 == result_fraction__492;
  assign eq_161743 = prod_bexp__46 == high_exp__92;
  assign eq_161744 = prod_fraction__33 == result_fraction__493;
  assign high_exp__385 = 8'hff;
  assign result_fraction__791 = 23'h00_0000;
  assign high_exp__386 = 8'hff;
  assign result_fraction__792 = 23'h00_0000;
  assign high_exp__158 = 8'hff;
  assign result_fraction__561 = 23'h00_0000;
  assign high_exp__159 = 8'hff;
  assign result_fraction__562 = 23'h00_0000;
  assign ne_161756 = x_fraction__187 != result_fraction__806;
  assign ne_161758 = prod_fraction__67 != result_fraction__807;
  assign eq_161759 = x_bexp__187 == high_exp__156;
  assign eq_161760 = x_fraction__187 == result_fraction__559;
  assign eq_161761 = prod_bexp__91 == high_exp__157;
  assign eq_161762 = prod_fraction__67 == result_fraction__560;
  assign high_exp__417 = 8'hff;
  assign result_fraction__824 = 23'h00_0000;
  assign high_exp__418 = 8'hff;
  assign result_fraction__825 = 23'h00_0000;
  assign high_exp__222 = 8'hff;
  assign result_fraction__624 = 23'h00_0000;
  assign high_exp__223 = 8'hff;
  assign result_fraction__625 = 23'h00_0000;
  assign ne_161775 = x_fraction__331 != result_fraction__839;
  assign ne_161777 = prod_fraction__121 != result_fraction__840;
  assign eq_161778 = x_bexp__331 == high_exp__220;
  assign eq_161779 = x_fraction__331 == result_fraction__622;
  assign eq_161780 = prod_bexp__163 == high_exp__221;
  assign eq_161781 = prod_fraction__121 == result_fraction__623;
  assign high_exp__449 = 8'hff;
  assign result_fraction__857 = 23'h00_0000;
  assign high_exp__450 = 8'hff;
  assign result_fraction__858 = 23'h00_0000;
  assign high_exp__292 = 8'hff;
  assign result_fraction__695 = 23'h00_0000;
  assign high_exp__293 = 8'hff;
  assign result_fraction__696 = 23'h00_0000;
  assign ne_161794 = x_fraction__475 != result_fraction__872;
  assign ne_161796 = prod_fraction__175 != result_fraction__873;
  assign eq_161797 = x_bexp__475 == high_exp__290;
  assign eq_161798 = x_fraction__475 == result_fraction__693;
  assign eq_161799 = prod_bexp__235 == high_exp__291;
  assign eq_161800 = prod_fraction__175 == result_fraction__694;
  assign ne_161803 = x_fraction__22 != result_fraction__758;
  assign ne_161805 = prod_fraction__7 != result_fraction__759;
  assign eq_161806 = x_bexp__22 == high_exp__93;
  assign eq_161807 = x_fraction__22 == result_fraction__494;
  assign eq_161808 = prod_bexp__10 == high_exp__94;
  assign eq_161809 = prod_fraction__7 == result_fraction__495;
  assign result_exp__10 = exp__16[8:0];
  assign ne_161820 = x_fraction__188 != result_fraction__791;
  assign ne_161822 = prod_fraction__68 != result_fraction__792;
  assign eq_161823 = x_bexp__188 == high_exp__158;
  assign eq_161824 = x_fraction__188 == result_fraction__561;
  assign eq_161825 = prod_bexp__92 == high_exp__159;
  assign eq_161826 = prod_fraction__68 == result_fraction__562;
  assign ne_161835 = x_fraction__332 != result_fraction__824;
  assign ne_161837 = prod_fraction__122 != result_fraction__825;
  assign eq_161838 = x_bexp__332 == high_exp__222;
  assign eq_161839 = x_fraction__332 == result_fraction__624;
  assign eq_161840 = prod_bexp__164 == high_exp__223;
  assign eq_161841 = prod_fraction__122 == result_fraction__625;
  assign result_exp__140 = exp__196[8:0];
  assign ne_161852 = x_fraction__476 != result_fraction__857;
  assign ne_161854 = prod_fraction__176 != result_fraction__858;
  assign eq_161855 = x_bexp__476 == high_exp__292;
  assign eq_161856 = x_fraction__476 == result_fraction__695;
  assign eq_161857 = prod_bexp__236 == high_exp__293;
  assign eq_161858 = prod_fraction__176 == result_fraction__696;
  assign result_exp__200 = exp__278[8:0];
  assign result_exp__11 = result_exp__10 & {9{$signed(exp__16) > $signed(10'h000)}};
  assign wide_exponent__35 = wide_exponent__34[8:0] & {9{~wide_exponent__34[9]}};
  assign has_pos_inf__11 = ~(x_bexp__94 != high_exp__367 | ne_161738 | x_sign__24) | ~(prod_bexp__46 != high_exp__368 | ne_161740 | prod_sign__11);
  assign has_neg_inf__11 = eq_161741 & eq_161742 & x_sign__24 | eq_161743 & eq_161744 & prod_sign__11;
  assign wide_exponent__74 = wide_exponent__72[8:0] & {9{~wide_exponent__72[9]}};
  assign has_pos_inf__24 = ~(x_bexp__187 != high_exp__399 | ne_161756 | x_sign__47) | ~(prod_bexp__91 != high_exp__400 | ne_161758 | prod_sign__23);
  assign has_neg_inf__24 = eq_161759 & eq_161760 & x_sign__47 | eq_161761 & eq_161762 & prod_sign__23;
  assign high_exp__226 = 8'hff;
  assign result_fraction__627 = 23'h00_0000;
  assign result_fraction__626 = 23'h00_0000;
  assign result_exp__142 = result_exp__140 & {9{$signed(exp__196) > $signed(10'h000)}};
  assign wide_exponent__131 = wide_exponent__129[8:0] & {9{~wide_exponent__129[9]}};
  assign has_pos_inf__43 = ~(x_bexp__331 != high_exp__431 | ne_161775 | x_sign__83) | ~(prod_bexp__163 != high_exp__432 | ne_161777 | prod_sign__41);
  assign has_neg_inf__43 = eq_161778 & eq_161779 & x_sign__83 | eq_161780 & eq_161781 & prod_sign__41;
  assign high_exp__296 = 8'hff;
  assign result_fraction__698 = 23'h00_0000;
  assign result_fraction__697 = 23'h00_0000;
  assign result_exp__202 = result_exp__200 & {9{$signed(exp__278) > $signed(10'h000)}};
  assign wide_exponent__188 = wide_exponent__186[8:0] & {9{~wide_exponent__186[9]}};
  assign has_pos_inf__62 = ~(x_bexp__475 != high_exp__463 | ne_161794 | x_sign__119) | ~(prod_bexp__235 != high_exp__464 | ne_161796 | prod_sign__59);
  assign has_neg_inf__62 = eq_161797 & eq_161798 & x_sign__119 | eq_161799 & eq_161800 & prod_sign__59;
  assign wide_exponent__9 = wide_exponent__8[8:0] & {9{~wide_exponent__8[9]}};
  assign has_pos_inf__3 = ~(x_bexp__22 != high_exp__353 | ne_161803 | x_sign__6) | ~(prod_bexp__10 != high_exp__354 | ne_161805 | prod_sign__3);
  assign has_neg_inf__3 = eq_161806 & eq_161807 & x_sign__6 | eq_161808 & eq_161809 & prod_sign__3;
  assign wide_exponent__75 = wide_exponent__73[8:0] & {9{~wide_exponent__73[9]}};
  assign has_pos_inf__25 = ~(x_bexp__188 != high_exp__385 | ne_161820 | x_sign__48) | ~(prod_bexp__92 != high_exp__386 | ne_161822 | prod_sign__24);
  assign has_neg_inf__25 = eq_161823 & eq_161824 & x_sign__48 | eq_161825 & eq_161826 & prod_sign__24;
  assign wide_exponent__132 = wide_exponent__130[8:0] & {9{~wide_exponent__130[9]}};
  assign has_pos_inf__44 = ~(x_bexp__332 != high_exp__417 | ne_161835 | x_sign__84) | ~(prod_bexp__164 != high_exp__418 | ne_161837 | prod_sign__42);
  assign has_neg_inf__44 = eq_161838 & eq_161839 & x_sign__84 | eq_161840 & eq_161841 & prod_sign__42;
  assign is_result_nan__91 = x_bexp__334 == high_exp__226;
  assign ne_161937 = x_fraction__334 != result_fraction__627;
  assign wide_exponent__189 = wide_exponent__187[8:0] & {9{~wide_exponent__187[9]}};
  assign has_pos_inf__63 = ~(x_bexp__476 != high_exp__449 | ne_161852 | x_sign__120) | ~(prod_bexp__236 != high_exp__450 | ne_161854 | prod_sign__60);
  assign has_neg_inf__63 = eq_161855 & eq_161856 & x_sign__120 | eq_161857 & eq_161858 & prod_sign__60;
  assign is_result_nan__130 = x_bexp__478 == high_exp__296;
  assign ne_161951 = x_fraction__478 != result_fraction__698;
  assign and_reduce_161969 = &result_exp__11[7:0];
  assign is_result_nan__23 = eq_161741 & ne_161738 | eq_161743 & ne_161740 | has_pos_inf__11 & has_neg_inf__11;
  assign is_operand_inf__11 = eq_161741 & eq_161742 | eq_161743 & eq_161744;
  assign and_reduce_161975 = &wide_exponent__35[7:0];
  assign is_result_nan__50 = eq_161759 & ne_161756 | eq_161761 & ne_161758 | has_pos_inf__24 & has_neg_inf__24;
  assign is_operand_inf__24 = eq_161759 & eq_161760 | eq_161761 & eq_161762;
  assign and_reduce_161988 = &wide_exponent__74[7:0];
  assign is_result_nan__92 = is_result_nan__91 & ne_161937;
  assign has_inf_arg__47 = is_result_nan__91 & x_fraction__334 == result_fraction__626;
  assign and_reduce_161999 = &result_exp__142[7:0];
  assign is_result_nan__89 = eq_161778 & ne_161775 | eq_161780 & ne_161777 | has_pos_inf__43 & has_neg_inf__43;
  assign is_operand_inf__43 = eq_161778 & eq_161779 | eq_161780 & eq_161781;
  assign and_reduce_162005 = &wide_exponent__131[7:0];
  assign is_result_nan__131 = is_result_nan__130 & ne_161951;
  assign has_inf_arg__67 = is_result_nan__130 & x_fraction__478 == result_fraction__697;
  assign and_reduce_162016 = &result_exp__202[7:0];
  assign is_result_nan__128 = eq_161797 & ne_161794 | eq_161799 & ne_161796 | has_pos_inf__62 & has_neg_inf__62;
  assign is_operand_inf__62 = eq_161797 & eq_161798 | eq_161799 & eq_161800;
  assign and_reduce_162022 = &wide_exponent__188[7:0];
  assign is_result_nan__6 = eq_161806 & ne_161803 | eq_161808 & ne_161805 | has_pos_inf__3 & has_neg_inf__3;
  assign is_operand_inf__3 = eq_161806 & eq_161807 | eq_161808 & eq_161809;
  assign and_reduce_162029 = &wide_exponent__9[7:0];
  assign high_exp__97 = 8'hff;
  assign fraction_shift__370 = 3'h3;
  assign fraction_shift__235 = 3'h4;
  assign high_exp__95 = 8'hff;
  assign result_exp__38 = {8{is_result_nan__24}};
  assign is_result_nan__51 = eq_161823 & ne_161820 | eq_161825 & ne_161822 | has_pos_inf__25 & has_neg_inf__25;
  assign is_operand_inf__25 = eq_161823 & eq_161824 | eq_161825 & eq_161826;
  assign and_reduce_162043 = &wide_exponent__75[7:0];
  assign fraction_shift__388 = 3'h3;
  assign fraction_shift__270 = 3'h4;
  assign high_exp__160 = 8'hff;
  assign is_result_nan__90 = eq_161838 & ne_161835 | eq_161840 & ne_161837 | has_pos_inf__44 & has_neg_inf__44;
  assign is_operand_inf__44 = eq_161838 & eq_161839 | eq_161840 & eq_161841;
  assign and_reduce_162055 = &wide_exponent__132[7:0];
  assign high_exp__227 = 8'hff;
  assign fraction_shift__406 = 3'h3;
  assign fraction_shift__305 = 3'h4;
  assign high_exp__224 = 8'hff;
  assign result_exp__143 = {8{is_result_nan__91}};
  assign is_result_nan__129 = eq_161855 & ne_161852 | eq_161857 & ne_161854 | has_pos_inf__63 & has_neg_inf__63;
  assign is_operand_inf__63 = eq_161855 & eq_161856 | eq_161857 & eq_161858;
  assign and_reduce_162070 = &wide_exponent__189[7:0];
  assign high_exp__297 = 8'hff;
  assign fraction_shift__424 = 3'h3;
  assign fraction_shift__340 = 3'h4;
  assign high_exp__294 = 8'hff;
  assign result_exp__203 = {8{is_result_nan__130}};
  assign fraction_shift__371 = 3'h3;
  assign fraction_shift__236 = 3'h4;
  assign is_subnormal__4 = $signed(exp__16) <= $signed(10'h000);
  assign high_exp__96 = 8'hff;
  assign result_exp__12 = is_result_nan__79 | has_inf_arg__41 | result_exp__11[8] | and_reduce_161969 ? high_exp__97 : result_exp__11[7:0];
  assign fraction_shift__36 = rounding_carry__11 ? fraction_shift__235 : fraction_shift__370;
  assign result_sign__412 = 1'h0;
  assign result_exponent__12 = is_result_nan__23 | is_operand_inf__11 | wide_exponent__35[8] | and_reduce_161975 ? high_exp__95 : wide_exponent__35[7:0];
  assign result_sign__413 = 1'h0;
  assign fraction_shift__389 = 3'h3;
  assign fraction_shift__271 = 3'h4;
  assign high_exp__161 = 8'hff;
  assign fraction_shift__74 = rounding_carry__24 ? fraction_shift__270 : fraction_shift__388;
  assign result_sign__509 = 1'h0;
  assign result_exponent__24 = is_result_nan__50 | is_operand_inf__24 | wide_exponent__74[8] | and_reduce_161988 ? high_exp__160 : wide_exponent__74[7:0];
  assign fraction_shift__407 = 3'h3;
  assign fraction_shift__306 = 3'h4;
  assign is_subnormal__48 = $signed(exp__196) <= $signed(10'h000);
  assign high_exp__225 = 8'hff;
  assign result_exp__144 = is_result_nan__92 | has_inf_arg__47 | result_exp__142[8] | and_reduce_161999 ? high_exp__227 : result_exp__142[7:0];
  assign fraction_shift__131 = rounding_carry__43 ? fraction_shift__305 : fraction_shift__406;
  assign result_sign__604 = 1'h0;
  assign result_exponent__43 = is_result_nan__89 | is_operand_inf__43 | wide_exponent__131[8] | and_reduce_162005 ? high_exp__224 : wide_exponent__131[7:0];
  assign result_sign__605 = 1'h0;
  assign fraction_shift__425 = 3'h3;
  assign fraction_shift__341 = 3'h4;
  assign is_subnormal__68 = $signed(exp__278) <= $signed(10'h000);
  assign high_exp__295 = 8'hff;
  assign result_exp__204 = is_result_nan__131 | has_inf_arg__67 | result_exp__202[8] | and_reduce_162016 ? high_exp__297 : result_exp__202[7:0];
  assign fraction_shift__188 = rounding_carry__62 ? fraction_shift__340 : fraction_shift__424;
  assign result_sign__710 = 1'h0;
  assign result_exponent__62 = is_result_nan__128 | is_operand_inf__62 | wide_exponent__188[8] | and_reduce_162022 ? high_exp__294 : wide_exponent__188[7:0];
  assign result_sign__711 = 1'h0;
  assign fraction_shift__9 = rounding_carry__3 ? fraction_shift__236 : fraction_shift__371;
  assign result_sign__414 = 1'h0;
  assign result_exponent__3 = is_result_nan__6 | is_operand_inf__3 | wide_exponent__9[8] | and_reduce_162029 ? high_exp__96 : wide_exponent__9[7:0];
  assign result_sign__415 = 1'h0;
  assign shrl_162134 = rounded_fraction__11 >> fraction_shift__36;
  assign fraction_shift__75 = rounding_carry__25 ? fraction_shift__271 : fraction_shift__389;
  assign result_sign__510 = 1'h0;
  assign result_exponent__25 = is_result_nan__51 | is_operand_inf__25 | wide_exponent__75[8] | and_reduce_162043 ? high_exp__161 : wide_exponent__75[7:0];
  assign shrl_162142 = rounded_fraction__24 >> fraction_shift__74;
  assign fraction_shift__132 = rounding_carry__44 ? fraction_shift__306 : fraction_shift__407;
  assign result_sign__606 = 1'h0;
  assign result_exponent__44 = is_result_nan__90 | is_operand_inf__44 | wide_exponent__132[8] | and_reduce_162055 ? high_exp__225 : wide_exponent__132[7:0];
  assign result_sign__607 = 1'h0;
  assign shrl_162152 = rounded_fraction__43 >> fraction_shift__131;
  assign fraction_shift__189 = rounding_carry__63 ? fraction_shift__341 : fraction_shift__425;
  assign result_sign__712 = 1'h0;
  assign result_exponent__63 = is_result_nan__129 | is_operand_inf__63 | wide_exponent__189[8] | and_reduce_162070 ? high_exp__295 : wide_exponent__189[7:0];
  assign result_sign__713 = 1'h0;
  assign shrl_162163 = rounded_fraction__62 >> fraction_shift__188;
  assign concat_162166 = {result_sign__711, ~result_exp__203};
  assign shrl_162167 = rounded_fraction__3 >> fraction_shift__9;
  assign result_fraction__69 = shrl_162134[22:0];
  assign sum__12 = {result_sign__412, result_exponent__12} + {result_sign__413, ~result_exp__38};
  assign shrl_162175 = rounded_fraction__25 >> fraction_shift__75;
  assign result_fraction__148 = shrl_162142[22:0];
  assign sum__26 = {result_sign__509, result_exponent__24} + concat_158878;
  assign shrl_162181 = rounded_fraction__44 >> fraction_shift__132;
  assign result_fraction__265 = shrl_162152[22:0];
  assign sum__45 = {result_sign__604, result_exponent__43} + {result_sign__605, ~result_exp__143};
  assign shrl_162189 = rounded_fraction__63 >> fraction_shift__189;
  assign concat_162193 = {result_sign__713, ~result_exp__204};
  assign result_fraction__382 = shrl_162163[22:0];
  assign sum__64 = {result_sign__710, result_exponent__62} + concat_162166;
  assign result_fraction__16 = shrl_162167[22:0];
  assign result_fraction__19 = fraction__35[22:0];
  assign sum__4 = {result_sign__414, result_exponent__3} + {result_sign__415, ~result_exp__12};
  assign result_fraction__70 = result_fraction__69 & {23{~(is_operand_inf__11 | wide_exponent__35[8] | and_reduce_161975 | ~((|wide_exponent__35[8:1]) | wide_exponent__35[0]))}};
  assign nan_fraction__86 = 23'h40_0000;
  assign result_fraction__149 = shrl_162175[22:0];
  assign sum__27 = {result_sign__510, result_exponent__25} + concat_158858;
  assign result_fraction__150 = result_fraction__148 & {23{~(is_operand_inf__24 | wide_exponent__74[8] | and_reduce_161988 | ~((|wide_exponent__74[8:1]) | wide_exponent__74[0]))}};
  assign nan_fraction__113 = 23'h40_0000;
  assign result_fraction__266 = shrl_162181[22:0];
  assign result_fraction__272 = fraction__428[22:0];
  assign sum__46 = {result_sign__606, result_exponent__44} + {result_sign__607, ~result_exp__144};
  assign result_fraction__267 = result_fraction__265 & {23{~(is_operand_inf__43 | wide_exponent__131[8] | and_reduce_162005 | ~((|wide_exponent__131[8:1]) | wide_exponent__131[0]))}};
  assign nan_fraction__140 = 23'h40_0000;
  assign result_fraction__383 = shrl_162189[22:0];
  assign result_fraction__389 = fraction__607[22:0];
  assign sum__65 = {result_sign__712, result_exponent__63} + concat_162193;
  assign result_fraction__384 = result_fraction__382 & {23{~(is_operand_inf__62 | wide_exponent__188[8] | and_reduce_162022 | ~((|wide_exponent__188[8:1]) | wide_exponent__188[0]))}};
  assign nan_fraction__169 = 23'h40_0000;
  assign result_fraction__17 = result_fraction__16 & {23{~(is_operand_inf__3 | wide_exponent__9[8] | and_reduce_162029 | ~((|wide_exponent__9[8:1]) | wide_exponent__9[0]))}};
  assign nan_fraction__87 = 23'h40_0000;
  assign result_fraction__20 = result_fraction__19 & {23{~(has_inf_arg__41 | result_exp__11[8] | and_reduce_161969 | is_subnormal__4)}};
  assign nan_fraction__88 = 23'h40_0000;
  assign result_fraction__71 = is_result_nan__23 ? nan_fraction__86 : result_fraction__70;
  assign result_fraction__473 = {is_result_nan__24, 22'h00_0000};
  assign prod_bexp__50 = sum__12[8] ? result_exp__38 : result_exponent__12;
  assign x_bexp__710 = 8'h00;
  assign result_fraction__151 = result_fraction__149 & {23{~(is_operand_inf__25 | wide_exponent__75[8] | and_reduce_162043 | ~((|wide_exponent__75[8:1]) | wide_exponent__75[0]))}};
  assign nan_fraction__114 = 23'h40_0000;
  assign result_fraction__152 = is_result_nan__50 ? nan_fraction__113 : result_fraction__150;
  assign prod_bexp__99 = sum__26[8] ? result_exp__132 : result_exponent__24;
  assign x_bexp__711 = 8'h00;
  assign result_fraction__268 = result_fraction__266 & {23{~(is_operand_inf__44 | wide_exponent__132[8] | and_reduce_162055 | ~((|wide_exponent__132[8:1]) | wide_exponent__132[0]))}};
  assign nan_fraction__141 = 23'h40_0000;
  assign result_fraction__274 = result_fraction__272 & {23{~(has_inf_arg__47 | result_exp__142[8] | and_reduce_161999 | is_subnormal__48)}};
  assign nan_fraction__142 = 23'h40_0000;
  assign result_fraction__269 = is_result_nan__89 ? nan_fraction__140 : result_fraction__267;
  assign result_fraction__474 = {is_result_nan__91, 22'h00_0000};
  assign prod_bexp__171 = sum__45[8] ? result_exp__143 : result_exponent__43;
  assign x_bexp__712 = 8'h00;
  assign result_fraction__385 = result_fraction__383 & {23{~(is_operand_inf__63 | wide_exponent__189[8] | and_reduce_162070 | ~((|wide_exponent__189[8:1]) | wide_exponent__189[0]))}};
  assign nan_fraction__170 = 23'h40_0000;
  assign result_fraction__391 = result_fraction__389 & {23{~(has_inf_arg__67 | result_exp__202[8] | and_reduce_162016 | is_subnormal__68)}};
  assign nan_fraction__171 = 23'h40_0000;
  assign result_fraction__386 = is_result_nan__128 ? nan_fraction__169 : result_fraction__384;
  assign result_fraction__475 = {is_result_nan__130, 22'h00_0000};
  assign prod_bexp__243 = sum__64[8] ? result_exp__203 : result_exponent__62;
  assign x_bexp__713 = 8'h00;
  assign result_fraction__18 = is_result_nan__6 ? nan_fraction__87 : result_fraction__17;
  assign result_fraction__21 = is_result_nan__79 ? nan_fraction__88 : result_fraction__20;
  assign prod_bexp__14 = sum__4[8] ? result_exp__12 : result_exponent__3;
  assign x_bexp__714 = 8'h00;
  assign fraction_is_zero__11 = add_161030 == 26'h000_0000 & xddend_y__11[2:0] == 3'h0;
  assign prod_fraction__36 = sum__12[8] ? result_fraction__473 : result_fraction__71;
  assign incremented_sum__82 = sum__12[7:0] + 8'h01;
  assign result_fraction__153 = is_result_nan__51 ? nan_fraction__114 : result_fraction__151;
  assign prod_bexp__100 = sum__27[8] ? result_exp__131 : result_exponent__25;
  assign x_bexp__715 = 8'h00;
  assign fraction_is_zero__24 = add_161033 == 26'h000_0000 & xddend_y__23[2:0] == 3'h0;
  assign prod_fraction__73 = sum__26[8] ? result_fraction__471 : result_fraction__152;
  assign incremented_sum__100 = sum__26[7:0] + 8'h01;
  assign result_fraction__270 = is_result_nan__90 ? nan_fraction__141 : result_fraction__268;
  assign result_fraction__276 = is_result_nan__92 ? nan_fraction__142 : result_fraction__274;
  assign prod_bexp__172 = sum__46[8] ? result_exp__144 : result_exponent__44;
  assign x_bexp__716 = 8'h00;
  assign fraction_is_zero__43 = add_161036 == 26'h000_0000 & xddend_y__41[2:0] == 3'h0;
  assign prod_fraction__127 = sum__45[8] ? result_fraction__474 : result_fraction__269;
  assign incremented_sum__118 = sum__45[7:0] + 8'h01;
  assign result_fraction__387 = is_result_nan__129 ? nan_fraction__170 : result_fraction__385;
  assign result_fraction__393 = is_result_nan__131 ? nan_fraction__171 : result_fraction__391;
  assign prod_bexp__244 = sum__65[8] ? result_exp__204 : result_exponent__63;
  assign x_bexp__717 = 8'h00;
  assign fraction_is_zero__62 = add_161039 == 26'h000_0000 & xddend_y__59[2:0] == 3'h0;
  assign prod_fraction__181 = sum__64[8] ? result_fraction__475 : result_fraction__386;
  assign incremented_sum__136 = sum__64[7:0] + 8'h01;
  assign fraction_is_zero__3 = add_161040 == 26'h000_0000 & xddend_y__3[2:0] == 3'h0;
  assign prod_fraction__10 = sum__4[8] ? result_fraction__21 : result_fraction__18;
  assign incremented_sum__83 = sum__4[7:0] + 8'h01;
  assign wide_y__24 = {2'h1, prod_fraction__36, 3'h0};
  assign x_bexpbs_difference__13 = sum__12[8] ? incremented_sum__82 : ~sum__12[7:0];
  assign fraction_is_zero__25 = add_161043 == 26'h000_0000 & xddend_y__24[2:0] == 3'h0;
  assign prod_fraction__74 = sum__27[8] ? result_fraction__251 : result_fraction__153;
  assign incremented_sum__101 = sum__27[7:0] + 8'h01;
  assign wide_y__51 = {2'h1, prod_fraction__73, 3'h0};
  assign x_bexpbs_difference__25 = sum__26[8] ? incremented_sum__100 : ~sum__26[7:0];
  assign fraction_is_zero__44 = add_161046 == 26'h000_0000 & xddend_y__42[2:0] == 3'h0;
  assign prod_fraction__128 = sum__46[8] ? result_fraction__276 : result_fraction__270;
  assign incremented_sum__119 = sum__46[7:0] + 8'h01;
  assign wide_y__89 = {2'h1, prod_fraction__127, 3'h0};
  assign x_bexpbs_difference__43 = sum__45[8] ? incremented_sum__118 : ~sum__45[7:0];
  assign fraction_is_zero__63 = add_161049 == 26'h000_0000 & xddend_y__60[2:0] == 3'h0;
  assign prod_fraction__182 = sum__65[8] ? result_fraction__393 : result_fraction__387;
  assign incremented_sum__137 = sum__65[7:0] + 8'h01;
  assign wide_y__127 = {2'h1, prod_fraction__181, 3'h0};
  assign x_bexpbs_difference__61 = sum__64[8] ? incremented_sum__136 : ~sum__64[7:0];
  assign wide_y__7 = {2'h1, prod_fraction__10, 3'h0};
  assign x_bexpbs_difference__4 = sum__4[8] ? incremented_sum__83 : ~sum__4[7:0];
  assign concat_162407 = {~(add_161030[25] | fraction_is_zero__11), add_161030[25], fraction_is_zero__11};
  assign x_bexp__102 = sum__12[8] ? result_exponent__12 : result_exp__38;
  assign x_bexp__718 = 8'h00;
  assign wide_y__25 = wide_y__24 & {28{prod_bexp__50 != x_bexp__710}};
  assign sub_162413 = 8'h1c - x_bexpbs_difference__13;
  assign wide_y__52 = {2'h1, prod_fraction__74, 3'h0};
  assign x_bexpbs_difference__26 = sum__27[8] ? incremented_sum__101 : ~sum__27[7:0];
  assign concat_162419 = {~(add_161033[25] | fraction_is_zero__24), add_161033[25], fraction_is_zero__24};
  assign x_bexp__203 = sum__26[8] ? result_exponent__24 : result_exp__132;
  assign x_bexp__719 = 8'h00;
  assign wide_y__53 = wide_y__51 & {28{prod_bexp__99 != x_bexp__711}};
  assign sub_162425 = 8'h1c - x_bexpbs_difference__25;
  assign wide_y__90 = {2'h1, prod_fraction__128, 3'h0};
  assign x_bexpbs_difference__44 = sum__46[8] ? incremented_sum__119 : ~sum__46[7:0];
  assign concat_162431 = {~(add_161036[25] | fraction_is_zero__43), add_161036[25], fraction_is_zero__43};
  assign x_bexp__347 = sum__45[8] ? result_exponent__43 : result_exp__143;
  assign x_bexp__720 = 8'h00;
  assign wide_y__91 = wide_y__89 & {28{prod_bexp__171 != x_bexp__712}};
  assign sub_162437 = 8'h1c - x_bexpbs_difference__43;
  assign wide_y__128 = {2'h1, prod_fraction__182, 3'h0};
  assign x_bexpbs_difference__62 = sum__65[8] ? incremented_sum__137 : ~sum__65[7:0];
  assign concat_162443 = {~(add_161039[25] | fraction_is_zero__62), add_161039[25], fraction_is_zero__62};
  assign x_bexp__491 = sum__64[8] ? result_exponent__62 : result_exp__203;
  assign x_bexp__721 = 8'h00;
  assign wide_y__129 = wide_y__127 & {28{prod_bexp__243 != x_bexp__713}};
  assign sub_162449 = 8'h1c - x_bexpbs_difference__61;
  assign concat_162450 = {~(add_161040[25] | fraction_is_zero__3), add_161040[25], fraction_is_zero__3};
  assign x_bexp__30 = sum__4[8] ? result_exponent__3 : result_exp__12;
  assign x_bexp__722 = 8'h00;
  assign wide_y__8 = wide_y__7 & {28{prod_bexp__14 != x_bexp__714}};
  assign sub_162456 = 8'h1c - x_bexpbs_difference__4;
  assign high_exp__480 = 8'hff;
  assign result_sign__57 = x_sign__24 & prod_sign__11 & concat_162407[0] | ~prod_sign__11 & concat_162407[1] | prod_sign__11 & concat_162407[2];
  assign x_fraction__102 = sum__12[8] ? result_fraction__71 : result_fraction__473;
  assign dropped__12 = sub_162413 >= 8'h1c ? 28'h000_0000 : wide_y__25 << sub_162413;
  assign concat_162465 = {~(add_161043[25] | fraction_is_zero__25), add_161043[25], fraction_is_zero__25};
  assign x_bexp__204 = sum__27[8] ? result_exponent__25 : result_exp__131;
  assign x_bexp__723 = 8'h00;
  assign wide_y__54 = wide_y__52 & {28{prod_bexp__100 != x_bexp__715}};
  assign sub_162471 = 8'h1c - x_bexpbs_difference__26;
  assign result_sign__122 = x_sign__47 & prod_sign__23 & concat_162419[0] | ~prod_sign__23 & concat_162419[1] | prod_sign__23 & concat_162419[2];
  assign x_fraction__203 = sum__26[8] ? result_fraction__152 : result_fraction__471;
  assign dropped__26 = sub_162425 >= 8'h1c ? 28'h000_0000 : wide_y__53 << sub_162425;
  assign concat_162479 = {~(add_161046[25] | fraction_is_zero__44), add_161046[25], fraction_is_zero__44};
  assign x_bexp__348 = sum__46[8] ? result_exponent__44 : result_exp__144;
  assign x_bexp__724 = 8'h00;
  assign wide_y__92 = wide_y__90 & {28{prod_bexp__172 != x_bexp__716}};
  assign sub_162485 = 8'h1c - x_bexpbs_difference__44;
  assign high_exp__484 = 8'hff;
  assign result_sign__219 = x_sign__83 & prod_sign__41 & concat_162431[0] | ~prod_sign__41 & concat_162431[1] | prod_sign__41 & concat_162431[2];
  assign x_fraction__347 = sum__45[8] ? result_fraction__269 : result_fraction__474;
  assign dropped__45 = sub_162437 >= 8'h1c ? 28'h000_0000 : wide_y__91 << sub_162437;
  assign concat_162494 = {~(add_161049[25] | fraction_is_zero__63), add_161049[25], fraction_is_zero__63};
  assign x_bexp__492 = sum__65[8] ? result_exponent__63 : result_exp__204;
  assign x_bexp__725 = 8'h00;
  assign wide_y__130 = wide_y__128 & {28{prod_bexp__244 != x_bexp__717}};
  assign sub_162500 = 8'h1c - x_bexpbs_difference__62;
  assign high_exp__487 = 8'hff;
  assign result_sign__316 = x_sign__119 & prod_sign__59 & concat_162443[0] | ~prod_sign__59 & concat_162443[1] | prod_sign__59 & concat_162443[2];
  assign x_fraction__491 = sum__64[8] ? result_fraction__386 : result_fraction__475;
  assign dropped__64 = sub_162449 >= 8'h1c ? 28'h000_0000 : wide_y__129 << sub_162449;
  assign result_sign__13 = x_sign__6 & prod_sign__3 & concat_162450[0] | ~prod_sign__3 & concat_162450[1] | prod_sign__3 & concat_162450[2];
  assign x_fraction__30 = sum__4[8] ? result_fraction__18 : result_fraction__21;
  assign dropped__4 = sub_162456 >= 8'h1c ? 28'h000_0000 : wide_y__8 << sub_162456;
  assign result_sign__58 = is_operand_inf__11 ? ~has_pos_inf__11 : result_sign__57;
  assign wide_x__24 = {2'h1, x_fraction__102, 3'h0};
  assign result_sign__123 = x_sign__48 & prod_sign__24 & concat_162465[0] | ~prod_sign__24 & concat_162465[1] | prod_sign__24 & concat_162465[2];
  assign x_fraction__204 = sum__27[8] ? result_fraction__153 : result_fraction__251;
  assign dropped__27 = sub_162471 >= 8'h1c ? 28'h000_0000 : wide_y__54 << sub_162471;
  assign result_sign__124 = is_operand_inf__24 ? ~has_pos_inf__24 : result_sign__122;
  assign wide_x__51 = {2'h1, x_fraction__203, 3'h0};
  assign x_sign__86 = array_index_161206[31:31];
  assign result_sign__220 = x_sign__84 & prod_sign__42 & concat_162479[0] | ~prod_sign__42 & concat_162479[1] | prod_sign__42 & concat_162479[2];
  assign x_fraction__348 = sum__46[8] ? result_fraction__270 : result_fraction__276;
  assign dropped__46 = sub_162485 >= 8'h1c ? 28'h000_0000 : wide_y__92 << sub_162485;
  assign result_sign__221 = is_operand_inf__43 ? ~has_pos_inf__43 : result_sign__219;
  assign wide_x__89 = {2'h1, x_fraction__347, 3'h0};
  assign x_sign__122 = array_index_161220[31:31];
  assign result_sign__317 = x_sign__120 & prod_sign__60 & concat_162494[0] | ~prod_sign__60 & concat_162494[1] | prod_sign__60 & concat_162494[2];
  assign x_fraction__492 = sum__65[8] ? result_fraction__387 : result_fraction__393;
  assign dropped__65 = sub_162500 >= 8'h1c ? 28'h000_0000 : wide_y__130 << sub_162500;
  assign result_sign__318 = is_operand_inf__62 ? ~has_pos_inf__62 : result_sign__316;
  assign wide_x__127 = {2'h1, x_fraction__491, 3'h0};
  assign result_sign__14 = is_operand_inf__3 ? ~has_pos_inf__3 : result_sign__13;
  assign wide_x__7 = {2'h1, x_fraction__30, 3'h0};
  assign result_sign__61 = x_bexp__289 != high_exp__480 & x_sign__73;
  assign result_sign__59 = ~is_result_nan__23 & result_sign__58;
  assign wide_x__25 = wide_x__24 & {28{x_bexp__102 != x_bexp__718}};
  assign result_sign__125 = is_operand_inf__25 ? ~has_pos_inf__25 : result_sign__123;
  assign wide_x__52 = {2'h1, x_fraction__204, 3'h0};
  assign result_sign__126 = ~is_result_nan__50 & result_sign__124;
  assign wide_x__53 = wide_x__51 & {28{x_bexp__203 != x_bexp__719}};
  assign nand_162587 = ~(is_result_nan__91 & ne_161937);
  assign result_sign__226 = ~x_sign__86;
  assign result_sign__222 = is_operand_inf__44 ? ~has_pos_inf__44 : result_sign__220;
  assign wide_x__90 = {2'h1, x_fraction__348, 3'h0};
  assign result_sign__227 = x_bexp__334 != high_exp__484 & x_sign__86;
  assign result_sign__223 = ~is_result_nan__89 & result_sign__221;
  assign wide_x__91 = wide_x__89 & {28{x_bexp__347 != x_bexp__720}};
  assign nand_162600 = ~(is_result_nan__130 & ne_161951);
  assign result_sign__323 = ~x_sign__122;
  assign result_sign__319 = is_operand_inf__63 ? ~has_pos_inf__63 : result_sign__317;
  assign wide_x__128 = {2'h1, x_fraction__492, 3'h0};
  assign result_sign__324 = x_bexp__478 != high_exp__487 & x_sign__122;
  assign result_sign__320 = ~is_result_nan__128 & result_sign__318;
  assign wide_x__129 = wide_x__127 & {28{x_bexp__491 != x_bexp__721}};
  assign result_sign__15 = ~is_result_nan__6 & result_sign__14;
  assign wide_x__8 = wide_x__7 & {28{x_bexp__30 != x_bexp__722}};
  assign x_sign__26 = sum__12[8] ? result_sign__59 : result_sign__61;
  assign prod_sign__12 = sum__12[8] ? result_sign__61 : result_sign__59;
  assign neg_162619 = -wide_x__25;
  assign sticky__38 = {27'h000_0000, dropped__12[27:3] != 25'h000_0000};
  assign result_sign__127 = ~is_result_nan__51 & result_sign__125;
  assign wide_x__54 = wide_x__52 & {28{x_bexp__204 != x_bexp__723}};
  assign x_sign__51 = sum__26[8] ? result_sign__126 : result_sign__208;
  assign prod_sign__25 = sum__26[8] ? result_sign__208 : result_sign__126;
  assign neg_162628 = -wide_x__53;
  assign sticky__82 = {27'h000_0000, dropped__26[27:3] != 25'h000_0000};
  assign result_sign__228 = nand_162587 & result_sign__226;
  assign result_sign__224 = ~is_result_nan__90 & result_sign__222;
  assign wide_x__92 = wide_x__90 & {28{x_bexp__348 != x_bexp__724}};
  assign x_sign__87 = sum__45[8] ? result_sign__223 : result_sign__227;
  assign prod_sign__43 = sum__45[8] ? result_sign__227 : result_sign__223;
  assign neg_162638 = -wide_x__91;
  assign sticky__141 = {27'h000_0000, dropped__45[27:3] != 25'h000_0000};
  assign result_sign__325 = nand_162600 & result_sign__323;
  assign result_sign__321 = ~is_result_nan__129 & result_sign__319;
  assign wide_x__130 = wide_x__128 & {28{x_bexp__492 != x_bexp__725}};
  assign x_sign__123 = sum__64[8] ? result_sign__320 : result_sign__324;
  assign prod_sign__61 = sum__64[8] ? result_sign__324 : result_sign__320;
  assign neg_162648 = -wide_x__129;
  assign sticky__200 = {27'h000_0000, dropped__64[27:3] != 25'h000_0000};
  assign x_sign__8 = sum__4[8] ? result_sign__15 : result_sign__197;
  assign prod_sign__4 = sum__4[8] ? result_sign__197 : result_sign__15;
  assign neg_162653 = -wide_x__8;
  assign sticky__12 = {27'h000_0000, dropped__4[27:3] != 25'h000_0000};
  assign xddend_y__12 = (x_bexpbs_difference__13 >= 8'h1c ? 28'h000_0000 : wide_y__25 >> x_bexpbs_difference__13) | sticky__38;
  assign x_sign__52 = sum__27[8] ? result_sign__127 : result_sign__294;
  assign prod_sign__26 = sum__27[8] ? result_sign__294 : result_sign__127;
  assign neg_162662 = -wide_x__54;
  assign sticky__83 = {27'h000_0000, dropped__27[27:3] != 25'h000_0000};
  assign xddend_y__25 = (x_bexpbs_difference__25 >= 8'h1c ? 28'h000_0000 : wide_y__53 >> x_bexpbs_difference__25) | sticky__82;
  assign x_sign__88 = sum__46[8] ? result_sign__224 : result_sign__228;
  assign prod_sign__44 = sum__46[8] ? result_sign__228 : result_sign__224;
  assign neg_162671 = -wide_x__92;
  assign sticky__142 = {27'h000_0000, dropped__46[27:3] != 25'h000_0000};
  assign xddend_y__43 = (x_bexpbs_difference__43 >= 8'h1c ? 28'h000_0000 : wide_y__91 >> x_bexpbs_difference__43) | sticky__141;
  assign x_sign__124 = sum__65[8] ? result_sign__321 : result_sign__325;
  assign prod_sign__62 = sum__65[8] ? result_sign__325 : result_sign__321;
  assign neg_162680 = -wide_x__130;
  assign sticky__201 = {27'h000_0000, dropped__65[27:3] != 25'h000_0000};
  assign xddend_y__61 = (x_bexpbs_difference__61 >= 8'h1c ? 28'h000_0000 : wide_y__129 >> x_bexpbs_difference__61) | sticky__200;
  assign xddend_y__4 = (x_bexpbs_difference__4 >= 8'h1c ? 28'h000_0000 : wide_y__8 >> x_bexpbs_difference__4) | sticky__12;
  assign sel_162691 = x_sign__26 ^ prod_sign__12 ? neg_162619[27:3] : wide_x__25[27:3];
  assign result_sign__999 = 1'h0;
  assign xddend_y__26 = (x_bexpbs_difference__26 >= 8'h1c ? 28'h000_0000 : wide_y__54 >> x_bexpbs_difference__26) | sticky__83;
  assign sel_162698 = x_sign__51 ^ prod_sign__25 ? neg_162628[27:3] : wide_x__53[27:3];
  assign result_sign__1000 = 1'h0;
  assign xddend_y__44 = (x_bexpbs_difference__44 >= 8'h1c ? 28'h000_0000 : wide_y__92 >> x_bexpbs_difference__44) | sticky__142;
  assign sel_162705 = x_sign__87 ^ prod_sign__43 ? neg_162638[27:3] : wide_x__91[27:3];
  assign result_sign__1001 = 1'h0;
  assign xddend_y__62 = (x_bexpbs_difference__62 >= 8'h1c ? 28'h000_0000 : wide_y__130 >> x_bexpbs_difference__62) | sticky__201;
  assign sel_162712 = x_sign__123 ^ prod_sign__61 ? neg_162648[27:3] : wide_x__129[27:3];
  assign result_sign__1002 = 1'h0;
  assign sel_162715 = x_sign__8 ^ prod_sign__4 ? neg_162653[27:3] : wide_x__8[27:3];
  assign result_sign__1003 = 1'h0;
  assign sel_162720 = x_sign__52 ^ prod_sign__26 ? neg_162662[27:3] : wide_x__54[27:3];
  assign result_sign__1004 = 1'h0;
  assign sel_162725 = x_sign__88 ^ prod_sign__44 ? neg_162671[27:3] : wide_x__92[27:3];
  assign result_sign__1005 = 1'h0;
  assign sel_162730 = x_sign__124 ^ prod_sign__62 ? neg_162680[27:3] : wide_x__130[27:3];
  assign result_sign__1006 = 1'h0;
  assign add_162737 = {{1{sel_162691[24]}}, sel_162691} + {result_sign__999, xddend_y__12[27:3]};
  assign add_162740 = {{1{sel_162698[24]}}, sel_162698} + {result_sign__1000, xddend_y__25[27:3]};
  assign add_162743 = {{1{sel_162705[24]}}, sel_162705} + {result_sign__1001, xddend_y__43[27:3]};
  assign add_162746 = {{1{sel_162712[24]}}, sel_162712} + {result_sign__1002, xddend_y__61[27:3]};
  assign add_162747 = {{1{sel_162715[24]}}, sel_162715} + {result_sign__1003, xddend_y__4[27:3]};
  assign add_162750 = {{1{sel_162720[24]}}, sel_162720} + {result_sign__1004, xddend_y__26[27:3]};
  assign add_162753 = {{1{sel_162725[24]}}, sel_162725} + {result_sign__1005, xddend_y__44[27:3]};
  assign add_162756 = {{1{sel_162730[24]}}, sel_162730} + {result_sign__1006, xddend_y__62[27:3]};
  assign concat_162761 = {add_162737[24:0], xddend_y__12[2:0]};
  assign concat_162764 = {add_162740[24:0], xddend_y__25[2:0]};
  assign concat_162767 = {add_162743[24:0], xddend_y__43[2:0]};
  assign concat_162770 = {add_162746[24:0], xddend_y__61[2:0]};
  assign concat_162771 = {add_162747[24:0], xddend_y__4[2:0]};
  assign concat_162774 = {add_162750[24:0], xddend_y__26[2:0]};
  assign concat_162777 = {add_162753[24:0], xddend_y__44[2:0]};
  assign concat_162780 = {add_162756[24:0], xddend_y__62[2:0]};
  assign xbs_fraction__12 = add_162737[25] ? -concat_162761 : concat_162761;
  assign xbs_fraction__25 = add_162740[25] ? -concat_162764 : concat_162764;
  assign xbs_fraction__43 = add_162743[25] ? -concat_162767 : concat_162767;
  assign xbs_fraction__61 = add_162746[25] ? -concat_162770 : concat_162770;
  assign xbs_fraction__4 = add_162747[25] ? -concat_162771 : concat_162771;
  assign reverse_162796 = {xbs_fraction__12[0], xbs_fraction__12[1], xbs_fraction__12[2], xbs_fraction__12[3], xbs_fraction__12[4], xbs_fraction__12[5], xbs_fraction__12[6], xbs_fraction__12[7], xbs_fraction__12[8], xbs_fraction__12[9], xbs_fraction__12[10], xbs_fraction__12[11], xbs_fraction__12[12], xbs_fraction__12[13], xbs_fraction__12[14], xbs_fraction__12[15], xbs_fraction__12[16], xbs_fraction__12[17], xbs_fraction__12[18], xbs_fraction__12[19], xbs_fraction__12[20], xbs_fraction__12[21], xbs_fraction__12[22], xbs_fraction__12[23], xbs_fraction__12[24], xbs_fraction__12[25], xbs_fraction__12[26], xbs_fraction__12[27]};
  assign xbs_fraction__26 = add_162750[25] ? -concat_162774 : concat_162774;
  assign reverse_162798 = {xbs_fraction__25[0], xbs_fraction__25[1], xbs_fraction__25[2], xbs_fraction__25[3], xbs_fraction__25[4], xbs_fraction__25[5], xbs_fraction__25[6], xbs_fraction__25[7], xbs_fraction__25[8], xbs_fraction__25[9], xbs_fraction__25[10], xbs_fraction__25[11], xbs_fraction__25[12], xbs_fraction__25[13], xbs_fraction__25[14], xbs_fraction__25[15], xbs_fraction__25[16], xbs_fraction__25[17], xbs_fraction__25[18], xbs_fraction__25[19], xbs_fraction__25[20], xbs_fraction__25[21], xbs_fraction__25[22], xbs_fraction__25[23], xbs_fraction__25[24], xbs_fraction__25[25], xbs_fraction__25[26], xbs_fraction__25[27]};
  assign xbs_fraction__44 = add_162753[25] ? -concat_162777 : concat_162777;
  assign reverse_162800 = {xbs_fraction__43[0], xbs_fraction__43[1], xbs_fraction__43[2], xbs_fraction__43[3], xbs_fraction__43[4], xbs_fraction__43[5], xbs_fraction__43[6], xbs_fraction__43[7], xbs_fraction__43[8], xbs_fraction__43[9], xbs_fraction__43[10], xbs_fraction__43[11], xbs_fraction__43[12], xbs_fraction__43[13], xbs_fraction__43[14], xbs_fraction__43[15], xbs_fraction__43[16], xbs_fraction__43[17], xbs_fraction__43[18], xbs_fraction__43[19], xbs_fraction__43[20], xbs_fraction__43[21], xbs_fraction__43[22], xbs_fraction__43[23], xbs_fraction__43[24], xbs_fraction__43[25], xbs_fraction__43[26], xbs_fraction__43[27]};
  assign xbs_fraction__62 = add_162756[25] ? -concat_162780 : concat_162780;
  assign reverse_162802 = {xbs_fraction__61[0], xbs_fraction__61[1], xbs_fraction__61[2], xbs_fraction__61[3], xbs_fraction__61[4], xbs_fraction__61[5], xbs_fraction__61[6], xbs_fraction__61[7], xbs_fraction__61[8], xbs_fraction__61[9], xbs_fraction__61[10], xbs_fraction__61[11], xbs_fraction__61[12], xbs_fraction__61[13], xbs_fraction__61[14], xbs_fraction__61[15], xbs_fraction__61[16], xbs_fraction__61[17], xbs_fraction__61[18], xbs_fraction__61[19], xbs_fraction__61[20], xbs_fraction__61[21], xbs_fraction__61[22], xbs_fraction__61[23], xbs_fraction__61[24], xbs_fraction__61[25], xbs_fraction__61[26], xbs_fraction__61[27]};
  assign reverse_162803 = {xbs_fraction__4[0], xbs_fraction__4[1], xbs_fraction__4[2], xbs_fraction__4[3], xbs_fraction__4[4], xbs_fraction__4[5], xbs_fraction__4[6], xbs_fraction__4[7], xbs_fraction__4[8], xbs_fraction__4[9], xbs_fraction__4[10], xbs_fraction__4[11], xbs_fraction__4[12], xbs_fraction__4[13], xbs_fraction__4[14], xbs_fraction__4[15], xbs_fraction__4[16], xbs_fraction__4[17], xbs_fraction__4[18], xbs_fraction__4[19], xbs_fraction__4[20], xbs_fraction__4[21], xbs_fraction__4[22], xbs_fraction__4[23], xbs_fraction__4[24], xbs_fraction__4[25], xbs_fraction__4[26], xbs_fraction__4[27]};
  assign one_hot_162804 = {reverse_162796[27:0] == 28'h000_0000, reverse_162796[27] && reverse_162796[26:0] == 27'h000_0000, reverse_162796[26] && reverse_162796[25:0] == 26'h000_0000, reverse_162796[25] && reverse_162796[24:0] == 25'h000_0000, reverse_162796[24] && reverse_162796[23:0] == 24'h00_0000, reverse_162796[23] && reverse_162796[22:0] == 23'h00_0000, reverse_162796[22] && reverse_162796[21:0] == 22'h00_0000, reverse_162796[21] && reverse_162796[20:0] == 21'h00_0000, reverse_162796[20] && reverse_162796[19:0] == 20'h0_0000, reverse_162796[19] && reverse_162796[18:0] == 19'h0_0000, reverse_162796[18] && reverse_162796[17:0] == 18'h0_0000, reverse_162796[17] && reverse_162796[16:0] == 17'h0_0000, reverse_162796[16] && reverse_162796[15:0] == 16'h0000, reverse_162796[15] && reverse_162796[14:0] == 15'h0000, reverse_162796[14] && reverse_162796[13:0] == 14'h0000, reverse_162796[13] && reverse_162796[12:0] == 13'h0000, reverse_162796[12] && reverse_162796[11:0] == 12'h000, reverse_162796[11] && reverse_162796[10:0] == 11'h000, reverse_162796[10] && reverse_162796[9:0] == 10'h000, reverse_162796[9] && reverse_162796[8:0] == 9'h000, reverse_162796[8] && reverse_162796[7:0] == 8'h00, reverse_162796[7] && reverse_162796[6:0] == 7'h00, reverse_162796[6] && reverse_162796[5:0] == 6'h00, reverse_162796[5] && reverse_162796[4:0] == 5'h00, reverse_162796[4] && reverse_162796[3:0] == 4'h0, reverse_162796[3] && reverse_162796[2:0] == 3'h0, reverse_162796[2] && reverse_162796[1:0] == 2'h0, reverse_162796[1] && !reverse_162796[0], reverse_162796[0]};
  assign reverse_162805 = {xbs_fraction__26[0], xbs_fraction__26[1], xbs_fraction__26[2], xbs_fraction__26[3], xbs_fraction__26[4], xbs_fraction__26[5], xbs_fraction__26[6], xbs_fraction__26[7], xbs_fraction__26[8], xbs_fraction__26[9], xbs_fraction__26[10], xbs_fraction__26[11], xbs_fraction__26[12], xbs_fraction__26[13], xbs_fraction__26[14], xbs_fraction__26[15], xbs_fraction__26[16], xbs_fraction__26[17], xbs_fraction__26[18], xbs_fraction__26[19], xbs_fraction__26[20], xbs_fraction__26[21], xbs_fraction__26[22], xbs_fraction__26[23], xbs_fraction__26[24], xbs_fraction__26[25], xbs_fraction__26[26], xbs_fraction__26[27]};
  assign one_hot_162806 = {reverse_162798[27:0] == 28'h000_0000, reverse_162798[27] && reverse_162798[26:0] == 27'h000_0000, reverse_162798[26] && reverse_162798[25:0] == 26'h000_0000, reverse_162798[25] && reverse_162798[24:0] == 25'h000_0000, reverse_162798[24] && reverse_162798[23:0] == 24'h00_0000, reverse_162798[23] && reverse_162798[22:0] == 23'h00_0000, reverse_162798[22] && reverse_162798[21:0] == 22'h00_0000, reverse_162798[21] && reverse_162798[20:0] == 21'h00_0000, reverse_162798[20] && reverse_162798[19:0] == 20'h0_0000, reverse_162798[19] && reverse_162798[18:0] == 19'h0_0000, reverse_162798[18] && reverse_162798[17:0] == 18'h0_0000, reverse_162798[17] && reverse_162798[16:0] == 17'h0_0000, reverse_162798[16] && reverse_162798[15:0] == 16'h0000, reverse_162798[15] && reverse_162798[14:0] == 15'h0000, reverse_162798[14] && reverse_162798[13:0] == 14'h0000, reverse_162798[13] && reverse_162798[12:0] == 13'h0000, reverse_162798[12] && reverse_162798[11:0] == 12'h000, reverse_162798[11] && reverse_162798[10:0] == 11'h000, reverse_162798[10] && reverse_162798[9:0] == 10'h000, reverse_162798[9] && reverse_162798[8:0] == 9'h000, reverse_162798[8] && reverse_162798[7:0] == 8'h00, reverse_162798[7] && reverse_162798[6:0] == 7'h00, reverse_162798[6] && reverse_162798[5:0] == 6'h00, reverse_162798[5] && reverse_162798[4:0] == 5'h00, reverse_162798[4] && reverse_162798[3:0] == 4'h0, reverse_162798[3] && reverse_162798[2:0] == 3'h0, reverse_162798[2] && reverse_162798[1:0] == 2'h0, reverse_162798[1] && !reverse_162798[0], reverse_162798[0]};
  assign reverse_162807 = {xbs_fraction__44[0], xbs_fraction__44[1], xbs_fraction__44[2], xbs_fraction__44[3], xbs_fraction__44[4], xbs_fraction__44[5], xbs_fraction__44[6], xbs_fraction__44[7], xbs_fraction__44[8], xbs_fraction__44[9], xbs_fraction__44[10], xbs_fraction__44[11], xbs_fraction__44[12], xbs_fraction__44[13], xbs_fraction__44[14], xbs_fraction__44[15], xbs_fraction__44[16], xbs_fraction__44[17], xbs_fraction__44[18], xbs_fraction__44[19], xbs_fraction__44[20], xbs_fraction__44[21], xbs_fraction__44[22], xbs_fraction__44[23], xbs_fraction__44[24], xbs_fraction__44[25], xbs_fraction__44[26], xbs_fraction__44[27]};
  assign one_hot_162808 = {reverse_162800[27:0] == 28'h000_0000, reverse_162800[27] && reverse_162800[26:0] == 27'h000_0000, reverse_162800[26] && reverse_162800[25:0] == 26'h000_0000, reverse_162800[25] && reverse_162800[24:0] == 25'h000_0000, reverse_162800[24] && reverse_162800[23:0] == 24'h00_0000, reverse_162800[23] && reverse_162800[22:0] == 23'h00_0000, reverse_162800[22] && reverse_162800[21:0] == 22'h00_0000, reverse_162800[21] && reverse_162800[20:0] == 21'h00_0000, reverse_162800[20] && reverse_162800[19:0] == 20'h0_0000, reverse_162800[19] && reverse_162800[18:0] == 19'h0_0000, reverse_162800[18] && reverse_162800[17:0] == 18'h0_0000, reverse_162800[17] && reverse_162800[16:0] == 17'h0_0000, reverse_162800[16] && reverse_162800[15:0] == 16'h0000, reverse_162800[15] && reverse_162800[14:0] == 15'h0000, reverse_162800[14] && reverse_162800[13:0] == 14'h0000, reverse_162800[13] && reverse_162800[12:0] == 13'h0000, reverse_162800[12] && reverse_162800[11:0] == 12'h000, reverse_162800[11] && reverse_162800[10:0] == 11'h000, reverse_162800[10] && reverse_162800[9:0] == 10'h000, reverse_162800[9] && reverse_162800[8:0] == 9'h000, reverse_162800[8] && reverse_162800[7:0] == 8'h00, reverse_162800[7] && reverse_162800[6:0] == 7'h00, reverse_162800[6] && reverse_162800[5:0] == 6'h00, reverse_162800[5] && reverse_162800[4:0] == 5'h00, reverse_162800[4] && reverse_162800[3:0] == 4'h0, reverse_162800[3] && reverse_162800[2:0] == 3'h0, reverse_162800[2] && reverse_162800[1:0] == 2'h0, reverse_162800[1] && !reverse_162800[0], reverse_162800[0]};
  assign reverse_162809 = {xbs_fraction__62[0], xbs_fraction__62[1], xbs_fraction__62[2], xbs_fraction__62[3], xbs_fraction__62[4], xbs_fraction__62[5], xbs_fraction__62[6], xbs_fraction__62[7], xbs_fraction__62[8], xbs_fraction__62[9], xbs_fraction__62[10], xbs_fraction__62[11], xbs_fraction__62[12], xbs_fraction__62[13], xbs_fraction__62[14], xbs_fraction__62[15], xbs_fraction__62[16], xbs_fraction__62[17], xbs_fraction__62[18], xbs_fraction__62[19], xbs_fraction__62[20], xbs_fraction__62[21], xbs_fraction__62[22], xbs_fraction__62[23], xbs_fraction__62[24], xbs_fraction__62[25], xbs_fraction__62[26], xbs_fraction__62[27]};
  assign one_hot_162810 = {reverse_162802[27:0] == 28'h000_0000, reverse_162802[27] && reverse_162802[26:0] == 27'h000_0000, reverse_162802[26] && reverse_162802[25:0] == 26'h000_0000, reverse_162802[25] && reverse_162802[24:0] == 25'h000_0000, reverse_162802[24] && reverse_162802[23:0] == 24'h00_0000, reverse_162802[23] && reverse_162802[22:0] == 23'h00_0000, reverse_162802[22] && reverse_162802[21:0] == 22'h00_0000, reverse_162802[21] && reverse_162802[20:0] == 21'h00_0000, reverse_162802[20] && reverse_162802[19:0] == 20'h0_0000, reverse_162802[19] && reverse_162802[18:0] == 19'h0_0000, reverse_162802[18] && reverse_162802[17:0] == 18'h0_0000, reverse_162802[17] && reverse_162802[16:0] == 17'h0_0000, reverse_162802[16] && reverse_162802[15:0] == 16'h0000, reverse_162802[15] && reverse_162802[14:0] == 15'h0000, reverse_162802[14] && reverse_162802[13:0] == 14'h0000, reverse_162802[13] && reverse_162802[12:0] == 13'h0000, reverse_162802[12] && reverse_162802[11:0] == 12'h000, reverse_162802[11] && reverse_162802[10:0] == 11'h000, reverse_162802[10] && reverse_162802[9:0] == 10'h000, reverse_162802[9] && reverse_162802[8:0] == 9'h000, reverse_162802[8] && reverse_162802[7:0] == 8'h00, reverse_162802[7] && reverse_162802[6:0] == 7'h00, reverse_162802[6] && reverse_162802[5:0] == 6'h00, reverse_162802[5] && reverse_162802[4:0] == 5'h00, reverse_162802[4] && reverse_162802[3:0] == 4'h0, reverse_162802[3] && reverse_162802[2:0] == 3'h0, reverse_162802[2] && reverse_162802[1:0] == 2'h0, reverse_162802[1] && !reverse_162802[0], reverse_162802[0]};
  assign one_hot_162811 = {reverse_162803[27:0] == 28'h000_0000, reverse_162803[27] && reverse_162803[26:0] == 27'h000_0000, reverse_162803[26] && reverse_162803[25:0] == 26'h000_0000, reverse_162803[25] && reverse_162803[24:0] == 25'h000_0000, reverse_162803[24] && reverse_162803[23:0] == 24'h00_0000, reverse_162803[23] && reverse_162803[22:0] == 23'h00_0000, reverse_162803[22] && reverse_162803[21:0] == 22'h00_0000, reverse_162803[21] && reverse_162803[20:0] == 21'h00_0000, reverse_162803[20] && reverse_162803[19:0] == 20'h0_0000, reverse_162803[19] && reverse_162803[18:0] == 19'h0_0000, reverse_162803[18] && reverse_162803[17:0] == 18'h0_0000, reverse_162803[17] && reverse_162803[16:0] == 17'h0_0000, reverse_162803[16] && reverse_162803[15:0] == 16'h0000, reverse_162803[15] && reverse_162803[14:0] == 15'h0000, reverse_162803[14] && reverse_162803[13:0] == 14'h0000, reverse_162803[13] && reverse_162803[12:0] == 13'h0000, reverse_162803[12] && reverse_162803[11:0] == 12'h000, reverse_162803[11] && reverse_162803[10:0] == 11'h000, reverse_162803[10] && reverse_162803[9:0] == 10'h000, reverse_162803[9] && reverse_162803[8:0] == 9'h000, reverse_162803[8] && reverse_162803[7:0] == 8'h00, reverse_162803[7] && reverse_162803[6:0] == 7'h00, reverse_162803[6] && reverse_162803[5:0] == 6'h00, reverse_162803[5] && reverse_162803[4:0] == 5'h00, reverse_162803[4] && reverse_162803[3:0] == 4'h0, reverse_162803[3] && reverse_162803[2:0] == 3'h0, reverse_162803[2] && reverse_162803[1:0] == 2'h0, reverse_162803[1] && !reverse_162803[0], reverse_162803[0]};
  assign encode_162812 = {one_hot_162804[16] | one_hot_162804[17] | one_hot_162804[18] | one_hot_162804[19] | one_hot_162804[20] | one_hot_162804[21] | one_hot_162804[22] | one_hot_162804[23] | one_hot_162804[24] | one_hot_162804[25] | one_hot_162804[26] | one_hot_162804[27] | one_hot_162804[28], one_hot_162804[8] | one_hot_162804[9] | one_hot_162804[10] | one_hot_162804[11] | one_hot_162804[12] | one_hot_162804[13] | one_hot_162804[14] | one_hot_162804[15] | one_hot_162804[24] | one_hot_162804[25] | one_hot_162804[26] | one_hot_162804[27] | one_hot_162804[28], one_hot_162804[4] | one_hot_162804[5] | one_hot_162804[6] | one_hot_162804[7] | one_hot_162804[12] | one_hot_162804[13] | one_hot_162804[14] | one_hot_162804[15] | one_hot_162804[20] | one_hot_162804[21] | one_hot_162804[22] | one_hot_162804[23] | one_hot_162804[28], one_hot_162804[2] | one_hot_162804[3] | one_hot_162804[6] | one_hot_162804[7] | one_hot_162804[10] | one_hot_162804[11] | one_hot_162804[14] | one_hot_162804[15] | one_hot_162804[18] | one_hot_162804[19] | one_hot_162804[22] | one_hot_162804[23] | one_hot_162804[26] | one_hot_162804[27], one_hot_162804[1] | one_hot_162804[3] | one_hot_162804[5] | one_hot_162804[7] | one_hot_162804[9] | one_hot_162804[11] | one_hot_162804[13] | one_hot_162804[15] | one_hot_162804[17] | one_hot_162804[19] | one_hot_162804[21] | one_hot_162804[23] | one_hot_162804[25] | one_hot_162804[27]};
  assign one_hot_162813 = {reverse_162805[27:0] == 28'h000_0000, reverse_162805[27] && reverse_162805[26:0] == 27'h000_0000, reverse_162805[26] && reverse_162805[25:0] == 26'h000_0000, reverse_162805[25] && reverse_162805[24:0] == 25'h000_0000, reverse_162805[24] && reverse_162805[23:0] == 24'h00_0000, reverse_162805[23] && reverse_162805[22:0] == 23'h00_0000, reverse_162805[22] && reverse_162805[21:0] == 22'h00_0000, reverse_162805[21] && reverse_162805[20:0] == 21'h00_0000, reverse_162805[20] && reverse_162805[19:0] == 20'h0_0000, reverse_162805[19] && reverse_162805[18:0] == 19'h0_0000, reverse_162805[18] && reverse_162805[17:0] == 18'h0_0000, reverse_162805[17] && reverse_162805[16:0] == 17'h0_0000, reverse_162805[16] && reverse_162805[15:0] == 16'h0000, reverse_162805[15] && reverse_162805[14:0] == 15'h0000, reverse_162805[14] && reverse_162805[13:0] == 14'h0000, reverse_162805[13] && reverse_162805[12:0] == 13'h0000, reverse_162805[12] && reverse_162805[11:0] == 12'h000, reverse_162805[11] && reverse_162805[10:0] == 11'h000, reverse_162805[10] && reverse_162805[9:0] == 10'h000, reverse_162805[9] && reverse_162805[8:0] == 9'h000, reverse_162805[8] && reverse_162805[7:0] == 8'h00, reverse_162805[7] && reverse_162805[6:0] == 7'h00, reverse_162805[6] && reverse_162805[5:0] == 6'h00, reverse_162805[5] && reverse_162805[4:0] == 5'h00, reverse_162805[4] && reverse_162805[3:0] == 4'h0, reverse_162805[3] && reverse_162805[2:0] == 3'h0, reverse_162805[2] && reverse_162805[1:0] == 2'h0, reverse_162805[1] && !reverse_162805[0], reverse_162805[0]};
  assign encode_162814 = {one_hot_162806[16] | one_hot_162806[17] | one_hot_162806[18] | one_hot_162806[19] | one_hot_162806[20] | one_hot_162806[21] | one_hot_162806[22] | one_hot_162806[23] | one_hot_162806[24] | one_hot_162806[25] | one_hot_162806[26] | one_hot_162806[27] | one_hot_162806[28], one_hot_162806[8] | one_hot_162806[9] | one_hot_162806[10] | one_hot_162806[11] | one_hot_162806[12] | one_hot_162806[13] | one_hot_162806[14] | one_hot_162806[15] | one_hot_162806[24] | one_hot_162806[25] | one_hot_162806[26] | one_hot_162806[27] | one_hot_162806[28], one_hot_162806[4] | one_hot_162806[5] | one_hot_162806[6] | one_hot_162806[7] | one_hot_162806[12] | one_hot_162806[13] | one_hot_162806[14] | one_hot_162806[15] | one_hot_162806[20] | one_hot_162806[21] | one_hot_162806[22] | one_hot_162806[23] | one_hot_162806[28], one_hot_162806[2] | one_hot_162806[3] | one_hot_162806[6] | one_hot_162806[7] | one_hot_162806[10] | one_hot_162806[11] | one_hot_162806[14] | one_hot_162806[15] | one_hot_162806[18] | one_hot_162806[19] | one_hot_162806[22] | one_hot_162806[23] | one_hot_162806[26] | one_hot_162806[27], one_hot_162806[1] | one_hot_162806[3] | one_hot_162806[5] | one_hot_162806[7] | one_hot_162806[9] | one_hot_162806[11] | one_hot_162806[13] | one_hot_162806[15] | one_hot_162806[17] | one_hot_162806[19] | one_hot_162806[21] | one_hot_162806[23] | one_hot_162806[25] | one_hot_162806[27]};
  assign one_hot_162815 = {reverse_162807[27:0] == 28'h000_0000, reverse_162807[27] && reverse_162807[26:0] == 27'h000_0000, reverse_162807[26] && reverse_162807[25:0] == 26'h000_0000, reverse_162807[25] && reverse_162807[24:0] == 25'h000_0000, reverse_162807[24] && reverse_162807[23:0] == 24'h00_0000, reverse_162807[23] && reverse_162807[22:0] == 23'h00_0000, reverse_162807[22] && reverse_162807[21:0] == 22'h00_0000, reverse_162807[21] && reverse_162807[20:0] == 21'h00_0000, reverse_162807[20] && reverse_162807[19:0] == 20'h0_0000, reverse_162807[19] && reverse_162807[18:0] == 19'h0_0000, reverse_162807[18] && reverse_162807[17:0] == 18'h0_0000, reverse_162807[17] && reverse_162807[16:0] == 17'h0_0000, reverse_162807[16] && reverse_162807[15:0] == 16'h0000, reverse_162807[15] && reverse_162807[14:0] == 15'h0000, reverse_162807[14] && reverse_162807[13:0] == 14'h0000, reverse_162807[13] && reverse_162807[12:0] == 13'h0000, reverse_162807[12] && reverse_162807[11:0] == 12'h000, reverse_162807[11] && reverse_162807[10:0] == 11'h000, reverse_162807[10] && reverse_162807[9:0] == 10'h000, reverse_162807[9] && reverse_162807[8:0] == 9'h000, reverse_162807[8] && reverse_162807[7:0] == 8'h00, reverse_162807[7] && reverse_162807[6:0] == 7'h00, reverse_162807[6] && reverse_162807[5:0] == 6'h00, reverse_162807[5] && reverse_162807[4:0] == 5'h00, reverse_162807[4] && reverse_162807[3:0] == 4'h0, reverse_162807[3] && reverse_162807[2:0] == 3'h0, reverse_162807[2] && reverse_162807[1:0] == 2'h0, reverse_162807[1] && !reverse_162807[0], reverse_162807[0]};
  assign encode_162816 = {one_hot_162808[16] | one_hot_162808[17] | one_hot_162808[18] | one_hot_162808[19] | one_hot_162808[20] | one_hot_162808[21] | one_hot_162808[22] | one_hot_162808[23] | one_hot_162808[24] | one_hot_162808[25] | one_hot_162808[26] | one_hot_162808[27] | one_hot_162808[28], one_hot_162808[8] | one_hot_162808[9] | one_hot_162808[10] | one_hot_162808[11] | one_hot_162808[12] | one_hot_162808[13] | one_hot_162808[14] | one_hot_162808[15] | one_hot_162808[24] | one_hot_162808[25] | one_hot_162808[26] | one_hot_162808[27] | one_hot_162808[28], one_hot_162808[4] | one_hot_162808[5] | one_hot_162808[6] | one_hot_162808[7] | one_hot_162808[12] | one_hot_162808[13] | one_hot_162808[14] | one_hot_162808[15] | one_hot_162808[20] | one_hot_162808[21] | one_hot_162808[22] | one_hot_162808[23] | one_hot_162808[28], one_hot_162808[2] | one_hot_162808[3] | one_hot_162808[6] | one_hot_162808[7] | one_hot_162808[10] | one_hot_162808[11] | one_hot_162808[14] | one_hot_162808[15] | one_hot_162808[18] | one_hot_162808[19] | one_hot_162808[22] | one_hot_162808[23] | one_hot_162808[26] | one_hot_162808[27], one_hot_162808[1] | one_hot_162808[3] | one_hot_162808[5] | one_hot_162808[7] | one_hot_162808[9] | one_hot_162808[11] | one_hot_162808[13] | one_hot_162808[15] | one_hot_162808[17] | one_hot_162808[19] | one_hot_162808[21] | one_hot_162808[23] | one_hot_162808[25] | one_hot_162808[27]};
  assign one_hot_162817 = {reverse_162809[27:0] == 28'h000_0000, reverse_162809[27] && reverse_162809[26:0] == 27'h000_0000, reverse_162809[26] && reverse_162809[25:0] == 26'h000_0000, reverse_162809[25] && reverse_162809[24:0] == 25'h000_0000, reverse_162809[24] && reverse_162809[23:0] == 24'h00_0000, reverse_162809[23] && reverse_162809[22:0] == 23'h00_0000, reverse_162809[22] && reverse_162809[21:0] == 22'h00_0000, reverse_162809[21] && reverse_162809[20:0] == 21'h00_0000, reverse_162809[20] && reverse_162809[19:0] == 20'h0_0000, reverse_162809[19] && reverse_162809[18:0] == 19'h0_0000, reverse_162809[18] && reverse_162809[17:0] == 18'h0_0000, reverse_162809[17] && reverse_162809[16:0] == 17'h0_0000, reverse_162809[16] && reverse_162809[15:0] == 16'h0000, reverse_162809[15] && reverse_162809[14:0] == 15'h0000, reverse_162809[14] && reverse_162809[13:0] == 14'h0000, reverse_162809[13] && reverse_162809[12:0] == 13'h0000, reverse_162809[12] && reverse_162809[11:0] == 12'h000, reverse_162809[11] && reverse_162809[10:0] == 11'h000, reverse_162809[10] && reverse_162809[9:0] == 10'h000, reverse_162809[9] && reverse_162809[8:0] == 9'h000, reverse_162809[8] && reverse_162809[7:0] == 8'h00, reverse_162809[7] && reverse_162809[6:0] == 7'h00, reverse_162809[6] && reverse_162809[5:0] == 6'h00, reverse_162809[5] && reverse_162809[4:0] == 5'h00, reverse_162809[4] && reverse_162809[3:0] == 4'h0, reverse_162809[3] && reverse_162809[2:0] == 3'h0, reverse_162809[2] && reverse_162809[1:0] == 2'h0, reverse_162809[1] && !reverse_162809[0], reverse_162809[0]};
  assign encode_162818 = {one_hot_162810[16] | one_hot_162810[17] | one_hot_162810[18] | one_hot_162810[19] | one_hot_162810[20] | one_hot_162810[21] | one_hot_162810[22] | one_hot_162810[23] | one_hot_162810[24] | one_hot_162810[25] | one_hot_162810[26] | one_hot_162810[27] | one_hot_162810[28], one_hot_162810[8] | one_hot_162810[9] | one_hot_162810[10] | one_hot_162810[11] | one_hot_162810[12] | one_hot_162810[13] | one_hot_162810[14] | one_hot_162810[15] | one_hot_162810[24] | one_hot_162810[25] | one_hot_162810[26] | one_hot_162810[27] | one_hot_162810[28], one_hot_162810[4] | one_hot_162810[5] | one_hot_162810[6] | one_hot_162810[7] | one_hot_162810[12] | one_hot_162810[13] | one_hot_162810[14] | one_hot_162810[15] | one_hot_162810[20] | one_hot_162810[21] | one_hot_162810[22] | one_hot_162810[23] | one_hot_162810[28], one_hot_162810[2] | one_hot_162810[3] | one_hot_162810[6] | one_hot_162810[7] | one_hot_162810[10] | one_hot_162810[11] | one_hot_162810[14] | one_hot_162810[15] | one_hot_162810[18] | one_hot_162810[19] | one_hot_162810[22] | one_hot_162810[23] | one_hot_162810[26] | one_hot_162810[27], one_hot_162810[1] | one_hot_162810[3] | one_hot_162810[5] | one_hot_162810[7] | one_hot_162810[9] | one_hot_162810[11] | one_hot_162810[13] | one_hot_162810[15] | one_hot_162810[17] | one_hot_162810[19] | one_hot_162810[21] | one_hot_162810[23] | one_hot_162810[25] | one_hot_162810[27]};
  assign encode_162819 = {one_hot_162811[16] | one_hot_162811[17] | one_hot_162811[18] | one_hot_162811[19] | one_hot_162811[20] | one_hot_162811[21] | one_hot_162811[22] | one_hot_162811[23] | one_hot_162811[24] | one_hot_162811[25] | one_hot_162811[26] | one_hot_162811[27] | one_hot_162811[28], one_hot_162811[8] | one_hot_162811[9] | one_hot_162811[10] | one_hot_162811[11] | one_hot_162811[12] | one_hot_162811[13] | one_hot_162811[14] | one_hot_162811[15] | one_hot_162811[24] | one_hot_162811[25] | one_hot_162811[26] | one_hot_162811[27] | one_hot_162811[28], one_hot_162811[4] | one_hot_162811[5] | one_hot_162811[6] | one_hot_162811[7] | one_hot_162811[12] | one_hot_162811[13] | one_hot_162811[14] | one_hot_162811[15] | one_hot_162811[20] | one_hot_162811[21] | one_hot_162811[22] | one_hot_162811[23] | one_hot_162811[28], one_hot_162811[2] | one_hot_162811[3] | one_hot_162811[6] | one_hot_162811[7] | one_hot_162811[10] | one_hot_162811[11] | one_hot_162811[14] | one_hot_162811[15] | one_hot_162811[18] | one_hot_162811[19] | one_hot_162811[22] | one_hot_162811[23] | one_hot_162811[26] | one_hot_162811[27], one_hot_162811[1] | one_hot_162811[3] | one_hot_162811[5] | one_hot_162811[7] | one_hot_162811[9] | one_hot_162811[11] | one_hot_162811[13] | one_hot_162811[15] | one_hot_162811[17] | one_hot_162811[19] | one_hot_162811[21] | one_hot_162811[23] | one_hot_162811[25] | one_hot_162811[27]};
  assign encode_162821 = {one_hot_162813[16] | one_hot_162813[17] | one_hot_162813[18] | one_hot_162813[19] | one_hot_162813[20] | one_hot_162813[21] | one_hot_162813[22] | one_hot_162813[23] | one_hot_162813[24] | one_hot_162813[25] | one_hot_162813[26] | one_hot_162813[27] | one_hot_162813[28], one_hot_162813[8] | one_hot_162813[9] | one_hot_162813[10] | one_hot_162813[11] | one_hot_162813[12] | one_hot_162813[13] | one_hot_162813[14] | one_hot_162813[15] | one_hot_162813[24] | one_hot_162813[25] | one_hot_162813[26] | one_hot_162813[27] | one_hot_162813[28], one_hot_162813[4] | one_hot_162813[5] | one_hot_162813[6] | one_hot_162813[7] | one_hot_162813[12] | one_hot_162813[13] | one_hot_162813[14] | one_hot_162813[15] | one_hot_162813[20] | one_hot_162813[21] | one_hot_162813[22] | one_hot_162813[23] | one_hot_162813[28], one_hot_162813[2] | one_hot_162813[3] | one_hot_162813[6] | one_hot_162813[7] | one_hot_162813[10] | one_hot_162813[11] | one_hot_162813[14] | one_hot_162813[15] | one_hot_162813[18] | one_hot_162813[19] | one_hot_162813[22] | one_hot_162813[23] | one_hot_162813[26] | one_hot_162813[27], one_hot_162813[1] | one_hot_162813[3] | one_hot_162813[5] | one_hot_162813[7] | one_hot_162813[9] | one_hot_162813[11] | one_hot_162813[13] | one_hot_162813[15] | one_hot_162813[17] | one_hot_162813[19] | one_hot_162813[21] | one_hot_162813[23] | one_hot_162813[25] | one_hot_162813[27]};
  assign encode_162823 = {one_hot_162815[16] | one_hot_162815[17] | one_hot_162815[18] | one_hot_162815[19] | one_hot_162815[20] | one_hot_162815[21] | one_hot_162815[22] | one_hot_162815[23] | one_hot_162815[24] | one_hot_162815[25] | one_hot_162815[26] | one_hot_162815[27] | one_hot_162815[28], one_hot_162815[8] | one_hot_162815[9] | one_hot_162815[10] | one_hot_162815[11] | one_hot_162815[12] | one_hot_162815[13] | one_hot_162815[14] | one_hot_162815[15] | one_hot_162815[24] | one_hot_162815[25] | one_hot_162815[26] | one_hot_162815[27] | one_hot_162815[28], one_hot_162815[4] | one_hot_162815[5] | one_hot_162815[6] | one_hot_162815[7] | one_hot_162815[12] | one_hot_162815[13] | one_hot_162815[14] | one_hot_162815[15] | one_hot_162815[20] | one_hot_162815[21] | one_hot_162815[22] | one_hot_162815[23] | one_hot_162815[28], one_hot_162815[2] | one_hot_162815[3] | one_hot_162815[6] | one_hot_162815[7] | one_hot_162815[10] | one_hot_162815[11] | one_hot_162815[14] | one_hot_162815[15] | one_hot_162815[18] | one_hot_162815[19] | one_hot_162815[22] | one_hot_162815[23] | one_hot_162815[26] | one_hot_162815[27], one_hot_162815[1] | one_hot_162815[3] | one_hot_162815[5] | one_hot_162815[7] | one_hot_162815[9] | one_hot_162815[11] | one_hot_162815[13] | one_hot_162815[15] | one_hot_162815[17] | one_hot_162815[19] | one_hot_162815[21] | one_hot_162815[23] | one_hot_162815[25] | one_hot_162815[27]};
  assign encode_162825 = {one_hot_162817[16] | one_hot_162817[17] | one_hot_162817[18] | one_hot_162817[19] | one_hot_162817[20] | one_hot_162817[21] | one_hot_162817[22] | one_hot_162817[23] | one_hot_162817[24] | one_hot_162817[25] | one_hot_162817[26] | one_hot_162817[27] | one_hot_162817[28], one_hot_162817[8] | one_hot_162817[9] | one_hot_162817[10] | one_hot_162817[11] | one_hot_162817[12] | one_hot_162817[13] | one_hot_162817[14] | one_hot_162817[15] | one_hot_162817[24] | one_hot_162817[25] | one_hot_162817[26] | one_hot_162817[27] | one_hot_162817[28], one_hot_162817[4] | one_hot_162817[5] | one_hot_162817[6] | one_hot_162817[7] | one_hot_162817[12] | one_hot_162817[13] | one_hot_162817[14] | one_hot_162817[15] | one_hot_162817[20] | one_hot_162817[21] | one_hot_162817[22] | one_hot_162817[23] | one_hot_162817[28], one_hot_162817[2] | one_hot_162817[3] | one_hot_162817[6] | one_hot_162817[7] | one_hot_162817[10] | one_hot_162817[11] | one_hot_162817[14] | one_hot_162817[15] | one_hot_162817[18] | one_hot_162817[19] | one_hot_162817[22] | one_hot_162817[23] | one_hot_162817[26] | one_hot_162817[27], one_hot_162817[1] | one_hot_162817[3] | one_hot_162817[5] | one_hot_162817[7] | one_hot_162817[9] | one_hot_162817[11] | one_hot_162817[13] | one_hot_162817[15] | one_hot_162817[17] | one_hot_162817[19] | one_hot_162817[21] | one_hot_162817[23] | one_hot_162817[25] | one_hot_162817[27]};
  assign cancel__13 = |encode_162812[4:1];
  assign carry_bit__12 = xbs_fraction__12[27];
  assign result_fraction__496 = 23'h00_0000;
  assign cancel__26 = |encode_162814[4:1];
  assign carry_bit__26 = xbs_fraction__25[27];
  assign result_fraction__563 = 23'h00_0000;
  assign cancel__45 = |encode_162816[4:1];
  assign carry_bit__45 = xbs_fraction__43[27];
  assign result_fraction__628 = 23'h00_0000;
  assign cancel__64 = |encode_162818[4:1];
  assign carry_bit__64 = xbs_fraction__61[27];
  assign result_fraction__699 = 23'h00_0000;
  assign cancel__4 = |encode_162819[4:1];
  assign carry_bit__4 = xbs_fraction__4[27];
  assign result_fraction__497 = 23'h00_0000;
  assign leading_zeroes__12 = {result_fraction__496, encode_162812};
  assign cancel__27 = |encode_162821[4:1];
  assign carry_bit__27 = xbs_fraction__26[27];
  assign result_fraction__564 = 23'h00_0000;
  assign leading_zeroes__26 = {result_fraction__563, encode_162814};
  assign cancel__46 = |encode_162823[4:1];
  assign carry_bit__46 = xbs_fraction__44[27];
  assign result_fraction__629 = 23'h00_0000;
  assign leading_zeroes__45 = {result_fraction__628, encode_162816};
  assign cancel__65 = |encode_162825[4:1];
  assign carry_bit__65 = xbs_fraction__62[27];
  assign result_fraction__700 = 23'h00_0000;
  assign leading_zeroes__64 = {result_fraction__699, encode_162818};
  assign leading_zeroes__4 = {result_fraction__497, encode_162819};
  assign carry_fraction__24 = xbs_fraction__12[27:1];
  assign add_162891 = leading_zeroes__12 + 28'hfff_ffff;
  assign leading_zeroes__27 = {result_fraction__564, encode_162821};
  assign carry_fraction__51 = xbs_fraction__25[27:1];
  assign add_162904 = leading_zeroes__26 + 28'hfff_ffff;
  assign leading_zeroes__46 = {result_fraction__629, encode_162823};
  assign carry_fraction__89 = xbs_fraction__43[27:1];
  assign add_162917 = leading_zeroes__45 + 28'hfff_ffff;
  assign leading_zeroes__65 = {result_fraction__700, encode_162825};
  assign carry_fraction__127 = xbs_fraction__61[27:1];
  assign add_162930 = leading_zeroes__64 + 28'hfff_ffff;
  assign carry_fraction__7 = xbs_fraction__4[27:1];
  assign add_162937 = leading_zeroes__4 + 28'hfff_ffff;
  assign concat_162938 = {~(carry_bit__12 | cancel__13), ~(carry_bit__12 | ~cancel__13), ~(~carry_bit__12 | cancel__13)};
  assign carry_fraction__25 = carry_fraction__24 | {26'h000_0000, xbs_fraction__12[0]};
  assign cancel_fraction__12 = add_162891 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__12[26:0] << add_162891;
  assign carry_fraction__52 = xbs_fraction__26[27:1];
  assign add_162947 = leading_zeroes__27 + 28'hfff_ffff;
  assign concat_162948 = {~(carry_bit__26 | cancel__26), ~(carry_bit__26 | ~cancel__26), ~(~carry_bit__26 | cancel__26)};
  assign carry_fraction__53 = carry_fraction__51 | {26'h000_0000, xbs_fraction__25[0]};
  assign cancel_fraction__26 = add_162904 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__25[26:0] << add_162904;
  assign carry_fraction__90 = xbs_fraction__44[27:1];
  assign add_162957 = leading_zeroes__46 + 28'hfff_ffff;
  assign concat_162958 = {~(carry_bit__45 | cancel__45), ~(carry_bit__45 | ~cancel__45), ~(~carry_bit__45 | cancel__45)};
  assign carry_fraction__91 = carry_fraction__89 | {26'h000_0000, xbs_fraction__43[0]};
  assign cancel_fraction__45 = add_162917 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__43[26:0] << add_162917;
  assign carry_fraction__128 = xbs_fraction__62[27:1];
  assign add_162967 = leading_zeroes__65 + 28'hfff_ffff;
  assign concat_162968 = {~(carry_bit__64 | cancel__64), ~(carry_bit__64 | ~cancel__64), ~(~carry_bit__64 | cancel__64)};
  assign carry_fraction__129 = carry_fraction__127 | {26'h000_0000, xbs_fraction__61[0]};
  assign cancel_fraction__64 = add_162930 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__61[26:0] << add_162930;
  assign concat_162971 = {~(carry_bit__4 | cancel__4), ~(carry_bit__4 | ~cancel__4), ~(~carry_bit__4 | cancel__4)};
  assign carry_fraction__8 = carry_fraction__7 | {26'h000_0000, xbs_fraction__4[0]};
  assign cancel_fraction__4 = add_162937 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__4[26:0] << add_162937;
  assign shifted_fraction__12 = carry_fraction__25 & {27{concat_162938[0]}} | cancel_fraction__12 & {27{concat_162938[1]}} | xbs_fraction__12[26:0] & {27{concat_162938[2]}};
  assign concat_162975 = {~(carry_bit__27 | cancel__27), ~(carry_bit__27 | ~cancel__27), ~(~carry_bit__27 | cancel__27)};
  assign carry_fraction__54 = carry_fraction__52 | {26'h000_0000, xbs_fraction__26[0]};
  assign cancel_fraction__27 = add_162947 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__26[26:0] << add_162947;
  assign shifted_fraction__26 = carry_fraction__53 & {27{concat_162948[0]}} | cancel_fraction__26 & {27{concat_162948[1]}} | xbs_fraction__25[26:0] & {27{concat_162948[2]}};
  assign concat_162979 = {~(carry_bit__46 | cancel__46), ~(carry_bit__46 | ~cancel__46), ~(~carry_bit__46 | cancel__46)};
  assign carry_fraction__92 = carry_fraction__90 | {26'h000_0000, xbs_fraction__44[0]};
  assign cancel_fraction__46 = add_162957 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__44[26:0] << add_162957;
  assign shifted_fraction__45 = carry_fraction__91 & {27{concat_162958[0]}} | cancel_fraction__45 & {27{concat_162958[1]}} | xbs_fraction__43[26:0] & {27{concat_162958[2]}};
  assign concat_162983 = {~(carry_bit__65 | cancel__65), ~(carry_bit__65 | ~cancel__65), ~(~carry_bit__65 | cancel__65)};
  assign carry_fraction__130 = carry_fraction__128 | {26'h000_0000, xbs_fraction__62[0]};
  assign cancel_fraction__65 = add_162967 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__62[26:0] << add_162967;
  assign shifted_fraction__64 = carry_fraction__129 & {27{concat_162968[0]}} | cancel_fraction__64 & {27{concat_162968[1]}} | xbs_fraction__61[26:0] & {27{concat_162968[2]}};
  assign shifted_fraction__4 = carry_fraction__8 & {27{concat_162971[0]}} | cancel_fraction__4 & {27{concat_162971[1]}} | xbs_fraction__4[26:0] & {27{concat_162971[2]}};
  assign result_sign__1007 = 1'h0;
  assign shifted_fraction__27 = carry_fraction__54 & {27{concat_162975[0]}} | cancel_fraction__27 & {27{concat_162975[1]}} | xbs_fraction__26[26:0] & {27{concat_162975[2]}};
  assign result_sign__1008 = 1'h0;
  assign shifted_fraction__46 = carry_fraction__92 & {27{concat_162979[0]}} | cancel_fraction__46 & {27{concat_162979[1]}} | xbs_fraction__44[26:0] & {27{concat_162979[2]}};
  assign result_sign__1009 = 1'h0;
  assign shifted_fraction__65 = carry_fraction__130 & {27{concat_162983[0]}} | cancel_fraction__65 & {27{concat_162983[1]}} | xbs_fraction__62[26:0] & {27{concat_162983[2]}};
  assign result_sign__1010 = 1'h0;
  assign result_sign__1011 = 1'h0;
  assign normal_chunk__12 = shifted_fraction__12[2:0];
  assign fraction_shift__237 = 3'h4;
  assign half_way_chunk__12 = shifted_fraction__12[3:2];
  assign result_sign__1012 = 1'h0;
  assign normal_chunk__26 = shifted_fraction__26[2:0];
  assign fraction_shift__272 = 3'h4;
  assign half_way_chunk__26 = shifted_fraction__26[3:2];
  assign result_sign__1013 = 1'h0;
  assign normal_chunk__45 = shifted_fraction__45[2:0];
  assign fraction_shift__307 = 3'h4;
  assign half_way_chunk__45 = shifted_fraction__45[3:2];
  assign result_sign__1014 = 1'h0;
  assign normal_chunk__64 = shifted_fraction__64[2:0];
  assign fraction_shift__342 = 3'h4;
  assign half_way_chunk__64 = shifted_fraction__64[3:2];
  assign normal_chunk__4 = shifted_fraction__4[2:0];
  assign fraction_shift__238 = 3'h4;
  assign half_way_chunk__4 = shifted_fraction__4[3:2];
  assign result_sign__416 = 1'h0;
  assign add_163040 = {result_sign__1007, shifted_fraction__12[26:3]} + 25'h000_0001;
  assign normal_chunk__27 = shifted_fraction__27[2:0];
  assign fraction_shift__273 = 3'h4;
  assign half_way_chunk__27 = shifted_fraction__27[3:2];
  assign result_sign__511 = 1'h0;
  assign add_163050 = {result_sign__1008, shifted_fraction__26[26:3]} + 25'h000_0001;
  assign normal_chunk__46 = shifted_fraction__46[2:0];
  assign fraction_shift__308 = 3'h4;
  assign half_way_chunk__46 = shifted_fraction__46[3:2];
  assign result_sign__608 = 1'h0;
  assign add_163060 = {result_sign__1009, shifted_fraction__45[26:3]} + 25'h000_0001;
  assign normal_chunk__65 = shifted_fraction__65[2:0];
  assign fraction_shift__343 = 3'h4;
  assign half_way_chunk__65 = shifted_fraction__65[3:2];
  assign result_sign__714 = 1'h0;
  assign add_163070 = {result_sign__1010, shifted_fraction__64[26:3]} + 25'h000_0001;
  assign result_sign__417 = 1'h0;
  assign add_163074 = {result_sign__1011, shifted_fraction__4[26:3]} + 25'h000_0001;
  assign do_round_up__25 = normal_chunk__12 > fraction_shift__237 | half_way_chunk__12 == 2'h3;
  assign result_sign__512 = 1'h0;
  assign add_163081 = {result_sign__1012, shifted_fraction__27[26:3]} + 25'h000_0001;
  assign do_round_up__54 = normal_chunk__26 > fraction_shift__272 | half_way_chunk__26 == 2'h3;
  assign result_sign__609 = 1'h0;
  assign add_163088 = {result_sign__1013, shifted_fraction__46[26:3]} + 25'h000_0001;
  assign do_round_up__93 = normal_chunk__45 > fraction_shift__307 | half_way_chunk__45 == 2'h3;
  assign result_sign__715 = 1'h0;
  assign add_163095 = {result_sign__1014, shifted_fraction__65[26:3]} + 25'h000_0001;
  assign do_round_up__132 = normal_chunk__64 > fraction_shift__342 | half_way_chunk__64 == 2'h3;
  assign do_round_up__8 = normal_chunk__4 > fraction_shift__238 | half_way_chunk__4 == 2'h3;
  assign rounded_fraction__12 = do_round_up__25 ? {add_163040, normal_chunk__12} : {result_sign__416, shifted_fraction__12};
  assign do_round_up__55 = normal_chunk__27 > fraction_shift__273 | half_way_chunk__27 == 2'h3;
  assign rounded_fraction__26 = do_round_up__54 ? {add_163050, normal_chunk__26} : {result_sign__511, shifted_fraction__26};
  assign do_round_up__94 = normal_chunk__46 > fraction_shift__308 | half_way_chunk__46 == 2'h3;
  assign rounded_fraction__45 = do_round_up__93 ? {add_163060, normal_chunk__45} : {result_sign__608, shifted_fraction__45};
  assign do_round_up__133 = normal_chunk__65 > fraction_shift__343 | half_way_chunk__65 == 2'h3;
  assign rounded_fraction__64 = do_round_up__132 ? {add_163070, normal_chunk__64} : {result_sign__714, shifted_fraction__64};
  assign rounded_fraction__4 = do_round_up__8 ? {add_163074, normal_chunk__4} : {result_sign__417, shifted_fraction__4};
  assign result_sign__418 = 1'h0;
  assign x_bexp__580 = 8'h00;
  assign rounding_carry__12 = rounded_fraction__12[27];
  assign rounded_fraction__27 = do_round_up__55 ? {add_163081, normal_chunk__27} : {result_sign__512, shifted_fraction__27};
  assign result_sign__513 = 1'h0;
  assign x_bexp__598 = 8'h00;
  assign rounding_carry__26 = rounded_fraction__26[27];
  assign rounded_fraction__46 = do_round_up__94 ? {add_163088, normal_chunk__46} : {result_sign__609, shifted_fraction__46};
  assign result_sign__610 = 1'h0;
  assign x_bexp__616 = 8'h00;
  assign rounding_carry__45 = rounded_fraction__45[27];
  assign rounded_fraction__65 = do_round_up__133 ? {add_163095, normal_chunk__65} : {result_sign__715, shifted_fraction__65};
  assign result_sign__716 = 1'h0;
  assign x_bexp__634 = 8'h00;
  assign rounding_carry__64 = rounded_fraction__64[27];
  assign result_sign__419 = 1'h0;
  assign x_bexp__581 = 8'h00;
  assign rounding_carry__4 = rounded_fraction__4[27];
  assign result_sign__514 = 1'h0;
  assign x_bexp__599 = 8'h00;
  assign rounding_carry__27 = rounded_fraction__27[27];
  assign result_sign__611 = 1'h0;
  assign x_bexp__617 = 8'h00;
  assign rounding_carry__46 = rounded_fraction__46[27];
  assign result_sign__717 = 1'h0;
  assign x_bexp__635 = 8'h00;
  assign rounding_carry__65 = rounded_fraction__65[27];
  assign result_sign__420 = 1'h0;
  assign add_163154 = {result_sign__418, x_bexp__102} + {x_bexp__580, rounding_carry__12};
  assign result_sign__515 = 1'h0;
  assign add_163160 = {result_sign__513, x_bexp__203} + {x_bexp__598, rounding_carry__26};
  assign result_sign__612 = 1'h0;
  assign add_163166 = {result_sign__610, x_bexp__347} + {x_bexp__616, rounding_carry__45};
  assign result_sign__718 = 1'h0;
  assign add_163172 = {result_sign__716, x_bexp__491} + {x_bexp__634, rounding_carry__64};
  assign result_sign__421 = 1'h0;
  assign add_163176 = {result_sign__419, x_bexp__30} + {x_bexp__581, rounding_carry__4};
  assign result_sign__516 = 1'h0;
  assign add_163185 = {result_sign__514, x_bexp__204} + {x_bexp__599, rounding_carry__27};
  assign result_sign__613 = 1'h0;
  assign add_163194 = {result_sign__611, x_bexp__348} + {x_bexp__617, rounding_carry__46};
  assign result_sign__719 = 1'h0;
  assign add_163203 = {result_sign__717, x_bexp__492} + {x_bexp__635, rounding_carry__65};
  assign add_163216 = {result_sign__420, add_163154} + 10'h001;
  assign add_163224 = {result_sign__515, add_163160} + 10'h001;
  assign add_163232 = {result_sign__612, add_163166} + 10'h001;
  assign add_163240 = {result_sign__718, add_163172} + 10'h001;
  assign add_163243 = {result_sign__421, add_163176} + 10'h001;
  assign wide_exponent__36 = add_163216 - {5'h00, encode_162812};
  assign add_163248 = {result_sign__516, add_163185} + 10'h001;
  assign wide_exponent__76 = add_163224 - {5'h00, encode_162814};
  assign add_163253 = {result_sign__613, add_163194} + 10'h001;
  assign wide_exponent__133 = add_163232 - {5'h00, encode_162816};
  assign add_163258 = {result_sign__719, add_163203} + 10'h001;
  assign wide_exponent__190 = add_163240 - {5'h00, encode_162818};
  assign wide_exponent__10 = add_163243 - {5'h00, encode_162819};
  assign wide_exponent__37 = wide_exponent__36 & {10{add_162737 != 26'h000_0000 | xddend_y__12[2:0] != 3'h0}};
  assign wide_exponent__77 = add_163248 - {5'h00, encode_162821};
  assign wide_exponent__78 = wide_exponent__76 & {10{add_162740 != 26'h000_0000 | xddend_y__25[2:0] != 3'h0}};
  assign wide_exponent__134 = add_163253 - {5'h00, encode_162823};
  assign wide_exponent__135 = wide_exponent__133 & {10{add_162743 != 26'h000_0000 | xddend_y__43[2:0] != 3'h0}};
  assign wide_exponent__191 = add_163258 - {5'h00, encode_162825};
  assign wide_exponent__192 = wide_exponent__190 & {10{add_162746 != 26'h000_0000 | xddend_y__61[2:0] != 3'h0}};
  assign wide_exponent__11 = wide_exponent__10 & {10{add_162747 != 26'h000_0000 | xddend_y__4[2:0] != 3'h0}};
  assign high_exp__369 = 8'hff;
  assign result_fraction__775 = 23'h00_0000;
  assign high_exp__370 = 8'hff;
  assign result_fraction__776 = 23'h00_0000;
  assign high_exp__98 = 8'hff;
  assign result_fraction__498 = 23'h00_0000;
  assign high_exp__99 = 8'hff;
  assign result_fraction__499 = 23'h00_0000;
  assign wide_exponent__79 = wide_exponent__77 & {10{add_162750 != 26'h000_0000 | xddend_y__26[2:0] != 3'h0}};
  assign high_exp__401 = 8'hff;
  assign result_fraction__808 = 23'h00_0000;
  assign high_exp__402 = 8'hff;
  assign result_fraction__809 = 23'h00_0000;
  assign high_exp__162 = 8'hff;
  assign result_fraction__565 = 23'h00_0000;
  assign high_exp__163 = 8'hff;
  assign result_fraction__566 = 23'h00_0000;
  assign wide_exponent__136 = wide_exponent__134 & {10{add_162753 != 26'h000_0000 | xddend_y__44[2:0] != 3'h0}};
  assign high_exp__433 = 8'hff;
  assign result_fraction__841 = 23'h00_0000;
  assign high_exp__434 = 8'hff;
  assign result_fraction__842 = 23'h00_0000;
  assign high_exp__228 = 8'hff;
  assign result_fraction__630 = 23'h00_0000;
  assign high_exp__229 = 8'hff;
  assign result_fraction__631 = 23'h00_0000;
  assign wide_exponent__193 = wide_exponent__191 & {10{add_162756 != 26'h000_0000 | xddend_y__62[2:0] != 3'h0}};
  assign high_exp__465 = 8'hff;
  assign result_fraction__874 = 23'h00_0000;
  assign high_exp__466 = 8'hff;
  assign result_fraction__875 = 23'h00_0000;
  assign high_exp__298 = 8'hff;
  assign result_fraction__701 = 23'h00_0000;
  assign high_exp__299 = 8'hff;
  assign result_fraction__702 = 23'h00_0000;
  assign high_exp__355 = 8'hff;
  assign result_fraction__760 = 23'h00_0000;
  assign high_exp__356 = 8'hff;
  assign result_fraction__761 = 23'h00_0000;
  assign high_exp__100 = 8'hff;
  assign result_fraction__500 = 23'h00_0000;
  assign high_exp__101 = 8'hff;
  assign result_fraction__501 = 23'h00_0000;
  assign ne_163326 = x_fraction__102 != result_fraction__775;
  assign ne_163328 = prod_fraction__36 != result_fraction__776;
  assign eq_163329 = x_bexp__102 == high_exp__98;
  assign eq_163330 = x_fraction__102 == result_fraction__498;
  assign eq_163331 = prod_bexp__50 == high_exp__99;
  assign eq_163332 = prod_fraction__36 == result_fraction__499;
  assign high_exp__387 = 8'hff;
  assign result_fraction__793 = 23'h00_0000;
  assign high_exp__388 = 8'hff;
  assign result_fraction__794 = 23'h00_0000;
  assign high_exp__164 = 8'hff;
  assign result_fraction__567 = 23'h00_0000;
  assign high_exp__165 = 8'hff;
  assign result_fraction__568 = 23'h00_0000;
  assign ne_163344 = x_fraction__203 != result_fraction__808;
  assign ne_163346 = prod_fraction__73 != result_fraction__809;
  assign eq_163347 = x_bexp__203 == high_exp__162;
  assign eq_163348 = x_fraction__203 == result_fraction__565;
  assign eq_163349 = prod_bexp__99 == high_exp__163;
  assign eq_163350 = prod_fraction__73 == result_fraction__566;
  assign high_exp__419 = 8'hff;
  assign result_fraction__826 = 23'h00_0000;
  assign high_exp__420 = 8'hff;
  assign result_fraction__827 = 23'h00_0000;
  assign high_exp__230 = 8'hff;
  assign result_fraction__632 = 23'h00_0000;
  assign high_exp__231 = 8'hff;
  assign result_fraction__633 = 23'h00_0000;
  assign ne_163362 = x_fraction__347 != result_fraction__841;
  assign ne_163364 = prod_fraction__127 != result_fraction__842;
  assign eq_163365 = x_bexp__347 == high_exp__228;
  assign eq_163366 = x_fraction__347 == result_fraction__630;
  assign eq_163367 = prod_bexp__171 == high_exp__229;
  assign eq_163368 = prod_fraction__127 == result_fraction__631;
  assign high_exp__451 = 8'hff;
  assign result_fraction__859 = 23'h00_0000;
  assign high_exp__452 = 8'hff;
  assign result_fraction__860 = 23'h00_0000;
  assign high_exp__300 = 8'hff;
  assign result_fraction__703 = 23'h00_0000;
  assign high_exp__301 = 8'hff;
  assign result_fraction__704 = 23'h00_0000;
  assign ne_163380 = x_fraction__491 != result_fraction__874;
  assign ne_163382 = prod_fraction__181 != result_fraction__875;
  assign eq_163383 = x_bexp__491 == high_exp__298;
  assign eq_163384 = x_fraction__491 == result_fraction__701;
  assign eq_163385 = prod_bexp__243 == high_exp__299;
  assign eq_163386 = prod_fraction__181 == result_fraction__702;
  assign ne_163389 = x_fraction__30 != result_fraction__760;
  assign ne_163391 = prod_fraction__10 != result_fraction__761;
  assign eq_163392 = x_bexp__30 == high_exp__100;
  assign eq_163393 = x_fraction__30 == result_fraction__500;
  assign eq_163394 = prod_bexp__14 == high_exp__101;
  assign eq_163395 = prod_fraction__10 == result_fraction__501;
  assign ne_163404 = x_fraction__204 != result_fraction__793;
  assign ne_163406 = prod_fraction__74 != result_fraction__794;
  assign eq_163407 = x_bexp__204 == high_exp__164;
  assign eq_163408 = x_fraction__204 == result_fraction__567;
  assign eq_163409 = prod_bexp__100 == high_exp__165;
  assign eq_163410 = prod_fraction__74 == result_fraction__568;
  assign ne_163419 = x_fraction__348 != result_fraction__826;
  assign ne_163421 = prod_fraction__128 != result_fraction__827;
  assign eq_163422 = x_bexp__348 == high_exp__230;
  assign eq_163423 = x_fraction__348 == result_fraction__632;
  assign eq_163424 = prod_bexp__172 == high_exp__231;
  assign eq_163425 = prod_fraction__128 == result_fraction__633;
  assign ne_163434 = x_fraction__492 != result_fraction__859;
  assign ne_163436 = prod_fraction__182 != result_fraction__860;
  assign eq_163437 = x_bexp__492 == high_exp__300;
  assign eq_163438 = x_fraction__492 == result_fraction__703;
  assign eq_163439 = prod_bexp__244 == high_exp__301;
  assign eq_163440 = prod_fraction__182 == result_fraction__704;
  assign wide_exponent__38 = wide_exponent__37[8:0] & {9{~wide_exponent__37[9]}};
  assign has_pos_inf__12 = ~(x_bexp__102 != high_exp__369 | ne_163326 | x_sign__26) | ~(prod_bexp__50 != high_exp__370 | ne_163328 | prod_sign__12);
  assign has_neg_inf__12 = eq_163329 & eq_163330 & x_sign__26 | eq_163331 & eq_163332 & prod_sign__12;
  assign wide_exponent__80 = wide_exponent__78[8:0] & {9{~wide_exponent__78[9]}};
  assign has_pos_inf__26 = ~(x_bexp__203 != high_exp__401 | ne_163344 | x_sign__51) | ~(prod_bexp__99 != high_exp__402 | ne_163346 | prod_sign__25);
  assign has_neg_inf__26 = eq_163347 & eq_163348 & x_sign__51 | eq_163349 & eq_163350 & prod_sign__25;
  assign wide_exponent__137 = wide_exponent__135[8:0] & {9{~wide_exponent__135[9]}};
  assign has_pos_inf__45 = ~(x_bexp__347 != high_exp__433 | ne_163362 | x_sign__87) | ~(prod_bexp__171 != high_exp__434 | ne_163364 | prod_sign__43);
  assign has_neg_inf__45 = eq_163365 & eq_163366 & x_sign__87 | eq_163367 & eq_163368 & prod_sign__43;
  assign wide_exponent__194 = wide_exponent__192[8:0] & {9{~wide_exponent__192[9]}};
  assign has_pos_inf__64 = ~(x_bexp__491 != high_exp__465 | ne_163380 | x_sign__123) | ~(prod_bexp__243 != high_exp__466 | ne_163382 | prod_sign__61);
  assign has_neg_inf__64 = eq_163383 & eq_163384 & x_sign__123 | eq_163385 & eq_163386 & prod_sign__61;
  assign array_index_163484 = in_img_unflattened[4'ha];
  assign wide_exponent__12 = wide_exponent__11[8:0] & {9{~wide_exponent__11[9]}};
  assign has_pos_inf__4 = ~(x_bexp__30 != high_exp__355 | ne_163389 | x_sign__8) | ~(prod_bexp__14 != high_exp__356 | ne_163391 | prod_sign__4);
  assign has_neg_inf__4 = eq_163392 & eq_163393 & x_sign__8 | eq_163394 & eq_163395 & prod_sign__4;
  assign wide_exponent__81 = wide_exponent__79[8:0] & {9{~wide_exponent__79[9]}};
  assign has_pos_inf__27 = ~(x_bexp__204 != high_exp__387 | ne_163404 | x_sign__52) | ~(prod_bexp__100 != high_exp__388 | ne_163406 | prod_sign__26);
  assign has_neg_inf__27 = eq_163407 & eq_163408 & x_sign__52 | eq_163409 & eq_163410 & prod_sign__26;
  assign wide_exponent__138 = wide_exponent__136[8:0] & {9{~wide_exponent__136[9]}};
  assign has_pos_inf__46 = ~(x_bexp__348 != high_exp__419 | ne_163419 | x_sign__88) | ~(prod_bexp__172 != high_exp__420 | ne_163421 | prod_sign__44);
  assign has_neg_inf__46 = eq_163422 & eq_163423 & x_sign__88 | eq_163424 & eq_163425 & prod_sign__44;
  assign wide_exponent__195 = wide_exponent__193[8:0] & {9{~wide_exponent__193[9]}};
  assign has_pos_inf__65 = ~(x_bexp__492 != high_exp__451 | ne_163434 | x_sign__124) | ~(prod_bexp__244 != high_exp__452 | ne_163436 | prod_sign__62);
  assign has_neg_inf__65 = eq_163437 & eq_163438 & x_sign__124 | eq_163439 & eq_163440 & prod_sign__62;
  assign x_bexp__503 = array_index_163484[30:23];
  assign high_exp__303 = 8'hff;
  assign is_result_nan__25 = eq_163329 & ne_163326 | eq_163331 & ne_163328 | has_pos_inf__12 & has_neg_inf__12;
  assign is_operand_inf__12 = eq_163329 & eq_163330 | eq_163331 & eq_163332;
  assign and_reduce_163539 = &wide_exponent__38[7:0];
  assign is_result_nan__54 = eq_163347 & ne_163344 | eq_163349 & ne_163346 | has_pos_inf__26 & has_neg_inf__26;
  assign is_operand_inf__26 = eq_163347 & eq_163348 | eq_163349 & eq_163350;
  assign and_reduce_163552 = &wide_exponent__80[7:0];
  assign is_result_nan__93 = eq_163365 & ne_163362 | eq_163367 & ne_163364 | has_pos_inf__45 & has_neg_inf__45;
  assign is_operand_inf__45 = eq_163365 & eq_163366 | eq_163367 & eq_163368;
  assign and_reduce_163565 = &wide_exponent__137[7:0];
  assign is_result_nan__132 = eq_163383 & ne_163380 | eq_163385 & ne_163382 | has_pos_inf__64 & has_neg_inf__64;
  assign is_operand_inf__64 = eq_163383 & eq_163384 | eq_163385 & eq_163386;
  assign and_reduce_163578 = &wide_exponent__194[7:0];
  assign is_result_nan__134 = x_bexp__503 == high_exp__303;
  assign is_result_nan__8 = eq_163392 & ne_163389 | eq_163394 & ne_163391 | has_pos_inf__4 & has_neg_inf__4;
  assign is_operand_inf__4 = eq_163392 & eq_163393 | eq_163394 & eq_163395;
  assign and_reduce_163585 = &wide_exponent__12[7:0];
  assign fraction_shift__372 = 3'h3;
  assign fraction_shift__239 = 3'h4;
  assign high_exp__102 = 8'hff;
  assign is_result_nan__55 = eq_163407 & ne_163404 | eq_163409 & ne_163406 | has_pos_inf__27 & has_neg_inf__27;
  assign is_operand_inf__27 = eq_163407 & eq_163408 | eq_163409 & eq_163410;
  assign and_reduce_163596 = &wide_exponent__81[7:0];
  assign fraction_shift__390 = 3'h3;
  assign fraction_shift__274 = 3'h4;
  assign high_exp__166 = 8'hff;
  assign is_result_nan__94 = eq_163422 & ne_163419 | eq_163424 & ne_163421 | has_pos_inf__46 & has_neg_inf__46;
  assign is_operand_inf__46 = eq_163422 & eq_163423 | eq_163424 & eq_163425;
  assign and_reduce_163607 = &wide_exponent__138[7:0];
  assign fraction_shift__408 = 3'h3;
  assign fraction_shift__309 = 3'h4;
  assign high_exp__232 = 8'hff;
  assign is_result_nan__133 = eq_163437 & ne_163434 | eq_163439 & ne_163436 | has_pos_inf__65 & has_neg_inf__65;
  assign is_operand_inf__65 = eq_163437 & eq_163438 | eq_163439 & eq_163440;
  assign and_reduce_163618 = &wide_exponent__195[7:0];
  assign fraction_shift__426 = 3'h3;
  assign fraction_shift__344 = 3'h4;
  assign high_exp__302 = 8'hff;
  assign result_exp__209 = {8{is_result_nan__134}};
  assign fraction_shift__373 = 3'h3;
  assign fraction_shift__240 = 3'h4;
  assign high_exp__103 = 8'hff;
  assign fraction_shift__39 = rounding_carry__12 ? fraction_shift__239 : fraction_shift__372;
  assign result_sign__422 = 1'h0;
  assign result_exponent__13 = is_result_nan__25 | is_operand_inf__12 | wide_exponent__38[8] | and_reduce_163539 ? high_exp__102 : wide_exponent__38[7:0];
  assign fraction_shift__391 = 3'h3;
  assign fraction_shift__275 = 3'h4;
  assign high_exp__167 = 8'hff;
  assign fraction_shift__80 = rounding_carry__26 ? fraction_shift__274 : fraction_shift__390;
  assign result_sign__517 = 1'h0;
  assign result_exponent__26 = is_result_nan__54 | is_operand_inf__26 | wide_exponent__80[8] | and_reduce_163552 ? high_exp__166 : wide_exponent__80[7:0];
  assign fraction_shift__409 = 3'h3;
  assign fraction_shift__310 = 3'h4;
  assign high_exp__233 = 8'hff;
  assign fraction_shift__137 = rounding_carry__45 ? fraction_shift__309 : fraction_shift__408;
  assign result_sign__614 = 1'h0;
  assign result_exponent__45 = is_result_nan__93 | is_operand_inf__45 | wide_exponent__137[8] | and_reduce_163565 ? high_exp__232 : wide_exponent__137[7:0];
  assign fraction_shift__427 = 3'h3;
  assign fraction_shift__345 = 3'h4;
  assign high_exp__304 = 8'hff;
  assign fraction_shift__194 = rounding_carry__64 ? fraction_shift__344 : fraction_shift__426;
  assign result_sign__720 = 1'h0;
  assign result_exponent__64 = is_result_nan__132 | is_operand_inf__64 | wide_exponent__194[8] | and_reduce_163578 ? high_exp__302 : wide_exponent__194[7:0];
  assign result_sign__721 = 1'h0;
  assign fraction_shift__12 = rounding_carry__4 ? fraction_shift__240 : fraction_shift__373;
  assign result_sign__423 = 1'h0;
  assign result_exponent__4 = is_result_nan__8 | is_operand_inf__4 | wide_exponent__12[8] | and_reduce_163585 ? high_exp__103 : wide_exponent__12[7:0];
  assign shrl_163667 = rounded_fraction__12 >> fraction_shift__39;
  assign fraction_shift__81 = rounding_carry__27 ? fraction_shift__275 : fraction_shift__391;
  assign result_sign__518 = 1'h0;
  assign result_exponent__27 = is_result_nan__55 | is_operand_inf__27 | wide_exponent__81[8] | and_reduce_163596 ? high_exp__167 : wide_exponent__81[7:0];
  assign shrl_163674 = rounded_fraction__26 >> fraction_shift__80;
  assign fraction_shift__138 = rounding_carry__46 ? fraction_shift__310 : fraction_shift__409;
  assign result_sign__615 = 1'h0;
  assign result_exponent__46 = is_result_nan__94 | is_operand_inf__46 | wide_exponent__138[8] | and_reduce_163607 ? high_exp__233 : wide_exponent__138[7:0];
  assign shrl_163681 = rounded_fraction__45 >> fraction_shift__137;
  assign fraction_shift__195 = rounding_carry__65 ? fraction_shift__345 : fraction_shift__427;
  assign result_sign__722 = 1'h0;
  assign result_exponent__65 = is_result_nan__133 | is_operand_inf__65 | wide_exponent__195[8] | and_reduce_163618 ? high_exp__304 : wide_exponent__195[7:0];
  assign shrl_163688 = rounded_fraction__64 >> fraction_shift__194;
  assign concat_163691 = {result_sign__721, ~result_exp__209};
  assign shrl_163692 = rounded_fraction__4 >> fraction_shift__12;
  assign result_fraction__75 = shrl_163667[22:0];
  assign sum__13 = {result_sign__422, result_exponent__13} + concat_158878;
  assign shrl_163698 = rounded_fraction__27 >> fraction_shift__81;
  assign result_fraction__160 = shrl_163674[22:0];
  assign sum__28 = {result_sign__517, result_exponent__26} + concat_158884;
  assign shrl_163704 = rounded_fraction__46 >> fraction_shift__138;
  assign result_fraction__277 = shrl_163681[22:0];
  assign sum__47 = {result_sign__614, result_exponent__45} + concat_162166;
  assign shrl_163710 = rounded_fraction__65 >> fraction_shift__195;
  assign result_fraction__394 = shrl_163688[22:0];
  assign sum__66 = {result_sign__720, result_exponent__64} + concat_163691;
  assign result_fraction__22 = shrl_163692[22:0];
  assign sum__5 = {result_sign__423, result_exponent__4} + concat_158878;
  assign result_fraction__76 = result_fraction__75 & {23{~(is_operand_inf__12 | wide_exponent__38[8] | and_reduce_163539 | ~((|wide_exponent__38[8:1]) | wide_exponent__38[0]))}};
  assign nan_fraction__89 = 23'h40_0000;
  assign result_fraction__161 = shrl_163698[22:0];
  assign sum__29 = {result_sign__518, result_exponent__27} + concat_158884;
  assign result_fraction__162 = result_fraction__160 & {23{~(is_operand_inf__26 | wide_exponent__80[8] | and_reduce_163552 | ~((|wide_exponent__80[8:1]) | wide_exponent__80[0]))}};
  assign nan_fraction__115 = 23'h40_0000;
  assign result_fraction__278 = shrl_163704[22:0];
  assign sum__48 = {result_sign__615, result_exponent__46} + concat_162166;
  assign result_fraction__279 = result_fraction__277 & {23{~(is_operand_inf__45 | wide_exponent__137[8] | and_reduce_163565 | ~((|wide_exponent__137[8:1]) | wide_exponent__137[0]))}};
  assign nan_fraction__143 = 23'h40_0000;
  assign result_fraction__395 = shrl_163710[22:0];
  assign sum__67 = {result_sign__722, result_exponent__65} + concat_163691;
  assign result_fraction__396 = result_fraction__394 & {23{~(is_operand_inf__64 | wide_exponent__194[8] | and_reduce_163578 | ~((|wide_exponent__194[8:1]) | wide_exponent__194[0]))}};
  assign nan_fraction__172 = 23'h40_0000;
  assign result_fraction__23 = result_fraction__22 & {23{~(is_operand_inf__4 | wide_exponent__12[8] | and_reduce_163585 | ~((|wide_exponent__12[8:1]) | wide_exponent__12[0]))}};
  assign nan_fraction__90 = 23'h40_0000;
  assign result_fraction__77 = is_result_nan__25 ? nan_fraction__89 : result_fraction__76;
  assign prod_bexp__54 = sum__13[8] ? result_exp__132 : result_exponent__13;
  assign x_bexp__726 = 8'h00;
  assign result_fraction__163 = result_fraction__161 & {23{~(is_operand_inf__27 | wide_exponent__81[8] | and_reduce_163596 | ~((|wide_exponent__81[8:1]) | wide_exponent__81[0]))}};
  assign nan_fraction__116 = 23'h40_0000;
  assign result_fraction__164 = is_result_nan__54 ? nan_fraction__115 : result_fraction__162;
  assign prod_bexp__107 = sum__28[8] ? result_exp__192 : result_exponent__26;
  assign x_bexp__727 = 8'h00;
  assign result_fraction__280 = result_fraction__278 & {23{~(is_operand_inf__46 | wide_exponent__138[8] | and_reduce_163607 | ~((|wide_exponent__138[8:1]) | wide_exponent__138[0]))}};
  assign nan_fraction__144 = 23'h40_0000;
  assign result_fraction__281 = is_result_nan__93 ? nan_fraction__143 : result_fraction__279;
  assign prod_bexp__179 = sum__47[8] ? result_exp__203 : result_exponent__45;
  assign x_bexp__728 = 8'h00;
  assign result_fraction__397 = result_fraction__395 & {23{~(is_operand_inf__65 | wide_exponent__195[8] | and_reduce_163618 | ~((|wide_exponent__195[8:1]) | wide_exponent__195[0]))}};
  assign nan_fraction__173 = 23'h40_0000;
  assign result_fraction__398 = is_result_nan__132 ? nan_fraction__172 : result_fraction__396;
  assign result_fraction__476 = {is_result_nan__134, 22'h00_0000};
  assign prod_bexp__251 = sum__66[8] ? result_exp__209 : result_exponent__64;
  assign x_bexp__729 = 8'h00;
  assign result_fraction__24 = is_result_nan__8 ? nan_fraction__90 : result_fraction__23;
  assign prod_bexp__18 = sum__5[8] ? result_exp__132 : result_exponent__4;
  assign x_bexp__730 = 8'h00;
  assign fraction_is_zero__12 = add_162737 == 26'h000_0000 & xddend_y__12[2:0] == 3'h0;
  assign prod_fraction__39 = sum__13[8] ? result_fraction__471 : result_fraction__77;
  assign incremented_sum__84 = sum__13[7:0] + 8'h01;
  assign result_fraction__165 = is_result_nan__55 ? nan_fraction__116 : result_fraction__163;
  assign prod_bexp__108 = sum__29[8] ? result_exp__192 : result_exponent__27;
  assign x_bexp__731 = 8'h00;
  assign fraction_is_zero__26 = add_162740 == 26'h000_0000 & xddend_y__25[2:0] == 3'h0;
  assign prod_fraction__79 = sum__28[8] ? result_fraction__472 : result_fraction__164;
  assign incremented_sum__102 = sum__28[7:0] + 8'h01;
  assign result_fraction__282 = is_result_nan__94 ? nan_fraction__144 : result_fraction__280;
  assign prod_bexp__180 = sum__48[8] ? result_exp__203 : result_exponent__46;
  assign x_bexp__732 = 8'h00;
  assign fraction_is_zero__45 = add_162743 == 26'h000_0000 & xddend_y__43[2:0] == 3'h0;
  assign prod_fraction__133 = sum__47[8] ? result_fraction__475 : result_fraction__281;
  assign incremented_sum__120 = sum__47[7:0] + 8'h01;
  assign result_fraction__399 = is_result_nan__133 ? nan_fraction__173 : result_fraction__397;
  assign prod_bexp__252 = sum__67[8] ? result_exp__209 : result_exponent__65;
  assign x_bexp__733 = 8'h00;
  assign fraction_is_zero__64 = add_162746 == 26'h000_0000 & xddend_y__61[2:0] == 3'h0;
  assign prod_fraction__187 = sum__66[8] ? result_fraction__476 : result_fraction__398;
  assign incremented_sum__138 = sum__66[7:0] + 8'h01;
  assign fraction_is_zero__4 = add_162747 == 26'h000_0000 & xddend_y__4[2:0] == 3'h0;
  assign prod_fraction__13 = sum__5[8] ? result_fraction__471 : result_fraction__24;
  assign incremented_sum__85 = sum__5[7:0] + 8'h01;
  assign wide_y__26 = {2'h1, prod_fraction__39, 3'h0};
  assign x_bexpbs_difference__14 = sum__13[8] ? incremented_sum__84 : ~sum__13[7:0];
  assign fraction_is_zero__27 = add_162750 == 26'h000_0000 & xddend_y__26[2:0] == 3'h0;
  assign prod_fraction__80 = sum__29[8] ? result_fraction__472 : result_fraction__165;
  assign incremented_sum__103 = sum__29[7:0] + 8'h01;
  assign wide_y__55 = {2'h1, prod_fraction__79, 3'h0};
  assign x_bexpbs_difference__27 = sum__28[8] ? incremented_sum__102 : ~sum__28[7:0];
  assign fraction_is_zero__46 = add_162753 == 26'h000_0000 & xddend_y__44[2:0] == 3'h0;
  assign prod_fraction__134 = sum__48[8] ? result_fraction__475 : result_fraction__282;
  assign incremented_sum__121 = sum__48[7:0] + 8'h01;
  assign wide_y__93 = {2'h1, prod_fraction__133, 3'h0};
  assign x_bexpbs_difference__45 = sum__47[8] ? incremented_sum__120 : ~sum__47[7:0];
  assign fraction_is_zero__65 = add_162756 == 26'h000_0000 & xddend_y__62[2:0] == 3'h0;
  assign prod_fraction__188 = sum__67[8] ? result_fraction__476 : result_fraction__399;
  assign incremented_sum__139 = sum__67[7:0] + 8'h01;
  assign wide_y__131 = {2'h1, prod_fraction__187, 3'h0};
  assign x_bexpbs_difference__63 = sum__66[8] ? incremented_sum__138 : ~sum__66[7:0];
  assign wide_y__9 = {2'h1, prod_fraction__13, 3'h0};
  assign x_bexpbs_difference__5 = sum__5[8] ? incremented_sum__85 : ~sum__5[7:0];
  assign concat_163907 = {~(add_162737[25] | fraction_is_zero__12), add_162737[25], fraction_is_zero__12};
  assign x_bexp__110 = sum__13[8] ? result_exponent__13 : result_exp__132;
  assign x_bexp__734 = 8'h00;
  assign wide_y__27 = wide_y__26 & {28{prod_bexp__54 != x_bexp__726}};
  assign sub_163913 = 8'h1c - x_bexpbs_difference__14;
  assign wide_y__56 = {2'h1, prod_fraction__80, 3'h0};
  assign x_bexpbs_difference__28 = sum__29[8] ? incremented_sum__103 : ~sum__29[7:0];
  assign concat_163919 = {~(add_162740[25] | fraction_is_zero__26), add_162740[25], fraction_is_zero__26};
  assign x_bexp__219 = sum__28[8] ? result_exponent__26 : result_exp__192;
  assign x_bexp__735 = 8'h00;
  assign wide_y__57 = wide_y__55 & {28{prod_bexp__107 != x_bexp__727}};
  assign sub_163925 = 8'h1c - x_bexpbs_difference__27;
  assign wide_y__94 = {2'h1, prod_fraction__134, 3'h0};
  assign x_bexpbs_difference__46 = sum__48[8] ? incremented_sum__121 : ~sum__48[7:0];
  assign concat_163931 = {~(add_162743[25] | fraction_is_zero__45), add_162743[25], fraction_is_zero__45};
  assign x_bexp__363 = sum__47[8] ? result_exponent__45 : result_exp__203;
  assign x_bexp__736 = 8'h00;
  assign wide_y__95 = wide_y__93 & {28{prod_bexp__179 != x_bexp__728}};
  assign sub_163937 = 8'h1c - x_bexpbs_difference__45;
  assign wide_y__132 = {2'h1, prod_fraction__188, 3'h0};
  assign x_bexpbs_difference__64 = sum__67[8] ? incremented_sum__139 : ~sum__67[7:0];
  assign concat_163943 = {~(add_162746[25] | fraction_is_zero__64), add_162746[25], fraction_is_zero__64};
  assign x_bexp__507 = sum__66[8] ? result_exponent__64 : result_exp__209;
  assign x_bexp__737 = 8'h00;
  assign wide_y__133 = wide_y__131 & {28{prod_bexp__251 != x_bexp__729}};
  assign sub_163949 = 8'h1c - x_bexpbs_difference__63;
  assign concat_163950 = {~(add_162747[25] | fraction_is_zero__4), add_162747[25], fraction_is_zero__4};
  assign x_bexp__38 = sum__5[8] ? result_exponent__4 : result_exp__132;
  assign x_bexp__738 = 8'h00;
  assign wide_y__10 = wide_y__9 & {28{prod_bexp__18 != x_bexp__730}};
  assign sub_163956 = 8'h1c - x_bexpbs_difference__5;
  assign result_sign__62 = x_sign__26 & prod_sign__12 & concat_163907[0] | ~prod_sign__12 & concat_163907[1] | prod_sign__12 & concat_163907[2];
  assign x_fraction__110 = sum__13[8] ? result_fraction__77 : result_fraction__471;
  assign dropped__13 = sub_163913 >= 8'h1c ? 28'h000_0000 : wide_y__27 << sub_163913;
  assign concat_163964 = {~(add_162750[25] | fraction_is_zero__27), add_162750[25], fraction_is_zero__27};
  assign x_bexp__220 = sum__29[8] ? result_exponent__27 : result_exp__192;
  assign x_bexp__739 = 8'h00;
  assign wide_y__58 = wide_y__56 & {28{prod_bexp__108 != x_bexp__731}};
  assign sub_163970 = 8'h1c - x_bexpbs_difference__28;
  assign result_sign__132 = x_sign__51 & prod_sign__25 & concat_163919[0] | ~prod_sign__25 & concat_163919[1] | prod_sign__25 & concat_163919[2];
  assign x_fraction__219 = sum__28[8] ? result_fraction__164 : result_fraction__472;
  assign dropped__28 = sub_163925 >= 8'h1c ? 28'h000_0000 : wide_y__57 << sub_163925;
  assign concat_163978 = {~(add_162753[25] | fraction_is_zero__46), add_162753[25], fraction_is_zero__46};
  assign x_bexp__364 = sum__48[8] ? result_exponent__46 : result_exp__203;
  assign x_bexp__740 = 8'h00;
  assign wide_y__96 = wide_y__94 & {28{prod_bexp__180 != x_bexp__732}};
  assign sub_163984 = 8'h1c - x_bexpbs_difference__46;
  assign result_sign__229 = x_sign__87 & prod_sign__43 & concat_163931[0] | ~prod_sign__43 & concat_163931[1] | prod_sign__43 & concat_163931[2];
  assign x_fraction__363 = sum__47[8] ? result_fraction__281 : result_fraction__475;
  assign dropped__47 = sub_163937 >= 8'h1c ? 28'h000_0000 : wide_y__95 << sub_163937;
  assign concat_163992 = {~(add_162756[25] | fraction_is_zero__65), add_162756[25], fraction_is_zero__65};
  assign x_bexp__508 = sum__67[8] ? result_exponent__65 : result_exp__209;
  assign x_bexp__741 = 8'h00;
  assign wide_y__134 = wide_y__132 & {28{prod_bexp__252 != x_bexp__733}};
  assign sub_163998 = 8'h1c - x_bexpbs_difference__64;
  assign high_exp__488 = 8'hff;
  assign result_sign__326 = x_sign__123 & prod_sign__61 & concat_163943[0] | ~prod_sign__61 & concat_163943[1] | prod_sign__61 & concat_163943[2];
  assign x_fraction__507 = sum__66[8] ? result_fraction__398 : result_fraction__476;
  assign dropped__66 = sub_163949 >= 8'h1c ? 28'h000_0000 : wide_y__133 << sub_163949;
  assign result_sign__18 = x_sign__8 & prod_sign__4 & concat_163950[0] | ~prod_sign__4 & concat_163950[1] | prod_sign__4 & concat_163950[2];
  assign x_fraction__38 = sum__5[8] ? result_fraction__24 : result_fraction__471;
  assign dropped__5 = sub_163956 >= 8'h1c ? 28'h000_0000 : wide_y__10 << sub_163956;
  assign result_sign__63 = is_operand_inf__12 ? ~has_pos_inf__12 : result_sign__62;
  assign wide_x__26 = {2'h1, x_fraction__110, 3'h0};
  assign result_sign__133 = x_sign__52 & prod_sign__26 & concat_163964[0] | ~prod_sign__26 & concat_163964[1] | prod_sign__26 & concat_163964[2];
  assign x_fraction__220 = sum__29[8] ? result_fraction__165 : result_fraction__472;
  assign dropped__29 = sub_163970 >= 8'h1c ? 28'h000_0000 : wide_y__58 << sub_163970;
  assign result_sign__134 = is_operand_inf__26 ? ~has_pos_inf__26 : result_sign__132;
  assign wide_x__55 = {2'h1, x_fraction__219, 3'h0};
  assign result_sign__230 = x_sign__88 & prod_sign__44 & concat_163978[0] | ~prod_sign__44 & concat_163978[1] | prod_sign__44 & concat_163978[2];
  assign x_fraction__364 = sum__48[8] ? result_fraction__282 : result_fraction__475;
  assign dropped__48 = sub_163984 >= 8'h1c ? 28'h000_0000 : wide_y__96 << sub_163984;
  assign result_sign__231 = is_operand_inf__45 ? ~has_pos_inf__45 : result_sign__229;
  assign wide_x__93 = {2'h1, x_fraction__363, 3'h0};
  assign result_sign__327 = x_sign__124 & prod_sign__62 & concat_163992[0] | ~prod_sign__62 & concat_163992[1] | prod_sign__62 & concat_163992[2];
  assign x_fraction__508 = sum__67[8] ? result_fraction__399 : result_fraction__476;
  assign dropped__67 = sub_163998 >= 8'h1c ? 28'h000_0000 : wide_y__134 << sub_163998;
  assign x_sign__125 = array_index_163484[31:31];
  assign result_sign__328 = is_operand_inf__64 ? ~has_pos_inf__64 : result_sign__326;
  assign wide_x__131 = {2'h1, x_fraction__507, 3'h0};
  assign result_sign__19 = is_operand_inf__4 ? ~has_pos_inf__4 : result_sign__18;
  assign wide_x__9 = {2'h1, x_fraction__38, 3'h0};
  assign result_sign__64 = ~is_result_nan__25 & result_sign__63;
  assign wide_x__27 = wide_x__26 & {28{x_bexp__110 != x_bexp__734}};
  assign result_sign__135 = is_operand_inf__27 ? ~has_pos_inf__27 : result_sign__133;
  assign wide_x__56 = {2'h1, x_fraction__220, 3'h0};
  assign result_sign__136 = ~is_result_nan__54 & result_sign__134;
  assign wide_x__57 = wide_x__55 & {28{x_bexp__219 != x_bexp__735}};
  assign result_sign__232 = is_operand_inf__46 ? ~has_pos_inf__46 : result_sign__230;
  assign wide_x__94 = {2'h1, x_fraction__364, 3'h0};
  assign result_sign__233 = ~is_result_nan__93 & result_sign__231;
  assign wide_x__95 = wide_x__93 & {28{x_bexp__363 != x_bexp__736}};
  assign result_sign__329 = is_operand_inf__65 ? ~has_pos_inf__65 : result_sign__327;
  assign wide_x__132 = {2'h1, x_fraction__508, 3'h0};
  assign result_sign__334 = x_bexp__503 != high_exp__488 & x_sign__125;
  assign result_sign__330 = ~is_result_nan__132 & result_sign__328;
  assign wide_x__133 = wide_x__131 & {28{x_bexp__507 != x_bexp__737}};
  assign result_sign__20 = ~is_result_nan__8 & result_sign__19;
  assign wide_x__10 = wide_x__9 & {28{x_bexp__38 != x_bexp__738}};
  assign x_sign__28 = sum__13[8] ? result_sign__64 : result_sign__208;
  assign prod_sign__13 = sum__13[8] ? result_sign__208 : result_sign__64;
  assign neg_164108 = -wide_x__27;
  assign sticky__41 = {27'h000_0000, dropped__13[27:3] != 25'h000_0000};
  assign result_sign__137 = ~is_result_nan__55 & result_sign__135;
  assign wide_x__58 = wide_x__56 & {28{x_bexp__220 != x_bexp__739}};
  assign x_sign__55 = sum__28[8] ? result_sign__136 : result_sign__305;
  assign prod_sign__27 = sum__28[8] ? result_sign__305 : result_sign__136;
  assign neg_164117 = -wide_x__57;
  assign sticky__88 = {27'h000_0000, dropped__28[27:3] != 25'h000_0000};
  assign result_sign__234 = ~is_result_nan__94 & result_sign__232;
  assign wide_x__96 = wide_x__94 & {28{x_bexp__364 != x_bexp__740}};
  assign x_sign__91 = sum__47[8] ? result_sign__233 : result_sign__324;
  assign prod_sign__45 = sum__47[8] ? result_sign__324 : result_sign__233;
  assign neg_164126 = -wide_x__95;
  assign sticky__147 = {27'h000_0000, dropped__47[27:3] != 25'h000_0000};
  assign result_sign__331 = ~is_result_nan__133 & result_sign__329;
  assign wide_x__134 = wide_x__132 & {28{x_bexp__508 != x_bexp__741}};
  assign x_sign__127 = sum__66[8] ? result_sign__330 : result_sign__334;
  assign prod_sign__63 = sum__66[8] ? result_sign__334 : result_sign__330;
  assign neg_164135 = -wide_x__133;
  assign sticky__206 = {27'h000_0000, dropped__66[27:3] != 25'h000_0000};
  assign x_sign__10 = sum__5[8] ? result_sign__20 : result_sign__208;
  assign prod_sign__5 = sum__5[8] ? result_sign__208 : result_sign__20;
  assign neg_164140 = -wide_x__10;
  assign sticky__15 = {27'h000_0000, dropped__5[27:3] != 25'h000_0000};
  assign xddend_y__13 = (x_bexpbs_difference__14 >= 8'h1c ? 28'h000_0000 : wide_y__27 >> x_bexpbs_difference__14) | sticky__41;
  assign x_sign__56 = sum__29[8] ? result_sign__137 : result_sign__305;
  assign prod_sign__28 = sum__29[8] ? result_sign__305 : result_sign__137;
  assign neg_164149 = -wide_x__58;
  assign sticky__89 = {27'h000_0000, dropped__29[27:3] != 25'h000_0000};
  assign xddend_y__27 = (x_bexpbs_difference__27 >= 8'h1c ? 28'h000_0000 : wide_y__57 >> x_bexpbs_difference__27) | sticky__88;
  assign x_sign__92 = sum__48[8] ? result_sign__234 : result_sign__324;
  assign prod_sign__46 = sum__48[8] ? result_sign__324 : result_sign__234;
  assign neg_164158 = -wide_x__96;
  assign sticky__148 = {27'h000_0000, dropped__48[27:3] != 25'h000_0000};
  assign xddend_y__45 = (x_bexpbs_difference__45 >= 8'h1c ? 28'h000_0000 : wide_y__95 >> x_bexpbs_difference__45) | sticky__147;
  assign x_sign__128 = sum__67[8] ? result_sign__331 : result_sign__334;
  assign prod_sign__64 = sum__67[8] ? result_sign__334 : result_sign__331;
  assign neg_164167 = -wide_x__134;
  assign sticky__207 = {27'h000_0000, dropped__67[27:3] != 25'h000_0000};
  assign xddend_y__63 = (x_bexpbs_difference__63 >= 8'h1c ? 28'h000_0000 : wide_y__133 >> x_bexpbs_difference__63) | sticky__206;
  assign xddend_y__5 = (x_bexpbs_difference__5 >= 8'h1c ? 28'h000_0000 : wide_y__10 >> x_bexpbs_difference__5) | sticky__15;
  assign sel_164178 = x_sign__28 ^ prod_sign__13 ? neg_164108[27:3] : wide_x__27[27:3];
  assign result_sign__1015 = 1'h0;
  assign xddend_y__28 = (x_bexpbs_difference__28 >= 8'h1c ? 28'h000_0000 : wide_y__58 >> x_bexpbs_difference__28) | sticky__89;
  assign sel_164185 = x_sign__55 ^ prod_sign__27 ? neg_164117[27:3] : wide_x__57[27:3];
  assign result_sign__1016 = 1'h0;
  assign xddend_y__46 = (x_bexpbs_difference__46 >= 8'h1c ? 28'h000_0000 : wide_y__96 >> x_bexpbs_difference__46) | sticky__148;
  assign sel_164192 = x_sign__91 ^ prod_sign__45 ? neg_164126[27:3] : wide_x__95[27:3];
  assign result_sign__1017 = 1'h0;
  assign xddend_y__64 = (x_bexpbs_difference__64 >= 8'h1c ? 28'h000_0000 : wide_y__134 >> x_bexpbs_difference__64) | sticky__207;
  assign sel_164199 = x_sign__127 ^ prod_sign__63 ? neg_164135[27:3] : wide_x__133[27:3];
  assign result_sign__1018 = 1'h0;
  assign sel_164202 = x_sign__10 ^ prod_sign__5 ? neg_164140[27:3] : wide_x__10[27:3];
  assign result_sign__1019 = 1'h0;
  assign sel_164207 = x_sign__56 ^ prod_sign__28 ? neg_164149[27:3] : wide_x__58[27:3];
  assign result_sign__1020 = 1'h0;
  assign sel_164212 = x_sign__92 ^ prod_sign__46 ? neg_164158[27:3] : wide_x__96[27:3];
  assign result_sign__1021 = 1'h0;
  assign sel_164217 = x_sign__128 ^ prod_sign__64 ? neg_164167[27:3] : wide_x__134[27:3];
  assign result_sign__1022 = 1'h0;
  assign add_164224 = {{1{sel_164178[24]}}, sel_164178} + {result_sign__1015, xddend_y__13[27:3]};
  assign add_164227 = {{1{sel_164185[24]}}, sel_164185} + {result_sign__1016, xddend_y__27[27:3]};
  assign add_164230 = {{1{sel_164192[24]}}, sel_164192} + {result_sign__1017, xddend_y__45[27:3]};
  assign add_164233 = {{1{sel_164199[24]}}, sel_164199} + {result_sign__1018, xddend_y__63[27:3]};
  assign add_164234 = {{1{sel_164202[24]}}, sel_164202} + {result_sign__1019, xddend_y__5[27:3]};
  assign add_164237 = {{1{sel_164207[24]}}, sel_164207} + {result_sign__1020, xddend_y__28[27:3]};
  assign add_164240 = {{1{sel_164212[24]}}, sel_164212} + {result_sign__1021, xddend_y__46[27:3]};
  assign add_164243 = {{1{sel_164217[24]}}, sel_164217} + {result_sign__1022, xddend_y__64[27:3]};
  assign concat_164248 = {add_164224[24:0], xddend_y__13[2:0]};
  assign concat_164251 = {add_164227[24:0], xddend_y__27[2:0]};
  assign concat_164254 = {add_164230[24:0], xddend_y__45[2:0]};
  assign concat_164257 = {add_164233[24:0], xddend_y__63[2:0]};
  assign concat_164258 = {add_164234[24:0], xddend_y__5[2:0]};
  assign concat_164261 = {add_164237[24:0], xddend_y__28[2:0]};
  assign concat_164264 = {add_164240[24:0], xddend_y__46[2:0]};
  assign concat_164267 = {add_164243[24:0], xddend_y__64[2:0]};
  assign xbs_fraction__13 = add_164224[25] ? -concat_164248 : concat_164248;
  assign xbs_fraction__27 = add_164227[25] ? -concat_164251 : concat_164251;
  assign xbs_fraction__45 = add_164230[25] ? -concat_164254 : concat_164254;
  assign xbs_fraction__63 = add_164233[25] ? -concat_164257 : concat_164257;
  assign xbs_fraction__5 = add_164234[25] ? -concat_164258 : concat_164258;
  assign reverse_164283 = {xbs_fraction__13[0], xbs_fraction__13[1], xbs_fraction__13[2], xbs_fraction__13[3], xbs_fraction__13[4], xbs_fraction__13[5], xbs_fraction__13[6], xbs_fraction__13[7], xbs_fraction__13[8], xbs_fraction__13[9], xbs_fraction__13[10], xbs_fraction__13[11], xbs_fraction__13[12], xbs_fraction__13[13], xbs_fraction__13[14], xbs_fraction__13[15], xbs_fraction__13[16], xbs_fraction__13[17], xbs_fraction__13[18], xbs_fraction__13[19], xbs_fraction__13[20], xbs_fraction__13[21], xbs_fraction__13[22], xbs_fraction__13[23], xbs_fraction__13[24], xbs_fraction__13[25], xbs_fraction__13[26], xbs_fraction__13[27]};
  assign xbs_fraction__28 = add_164237[25] ? -concat_164261 : concat_164261;
  assign reverse_164285 = {xbs_fraction__27[0], xbs_fraction__27[1], xbs_fraction__27[2], xbs_fraction__27[3], xbs_fraction__27[4], xbs_fraction__27[5], xbs_fraction__27[6], xbs_fraction__27[7], xbs_fraction__27[8], xbs_fraction__27[9], xbs_fraction__27[10], xbs_fraction__27[11], xbs_fraction__27[12], xbs_fraction__27[13], xbs_fraction__27[14], xbs_fraction__27[15], xbs_fraction__27[16], xbs_fraction__27[17], xbs_fraction__27[18], xbs_fraction__27[19], xbs_fraction__27[20], xbs_fraction__27[21], xbs_fraction__27[22], xbs_fraction__27[23], xbs_fraction__27[24], xbs_fraction__27[25], xbs_fraction__27[26], xbs_fraction__27[27]};
  assign xbs_fraction__46 = add_164240[25] ? -concat_164264 : concat_164264;
  assign reverse_164287 = {xbs_fraction__45[0], xbs_fraction__45[1], xbs_fraction__45[2], xbs_fraction__45[3], xbs_fraction__45[4], xbs_fraction__45[5], xbs_fraction__45[6], xbs_fraction__45[7], xbs_fraction__45[8], xbs_fraction__45[9], xbs_fraction__45[10], xbs_fraction__45[11], xbs_fraction__45[12], xbs_fraction__45[13], xbs_fraction__45[14], xbs_fraction__45[15], xbs_fraction__45[16], xbs_fraction__45[17], xbs_fraction__45[18], xbs_fraction__45[19], xbs_fraction__45[20], xbs_fraction__45[21], xbs_fraction__45[22], xbs_fraction__45[23], xbs_fraction__45[24], xbs_fraction__45[25], xbs_fraction__45[26], xbs_fraction__45[27]};
  assign xbs_fraction__64 = add_164243[25] ? -concat_164267 : concat_164267;
  assign reverse_164289 = {xbs_fraction__63[0], xbs_fraction__63[1], xbs_fraction__63[2], xbs_fraction__63[3], xbs_fraction__63[4], xbs_fraction__63[5], xbs_fraction__63[6], xbs_fraction__63[7], xbs_fraction__63[8], xbs_fraction__63[9], xbs_fraction__63[10], xbs_fraction__63[11], xbs_fraction__63[12], xbs_fraction__63[13], xbs_fraction__63[14], xbs_fraction__63[15], xbs_fraction__63[16], xbs_fraction__63[17], xbs_fraction__63[18], xbs_fraction__63[19], xbs_fraction__63[20], xbs_fraction__63[21], xbs_fraction__63[22], xbs_fraction__63[23], xbs_fraction__63[24], xbs_fraction__63[25], xbs_fraction__63[26], xbs_fraction__63[27]};
  assign reverse_164290 = {xbs_fraction__5[0], xbs_fraction__5[1], xbs_fraction__5[2], xbs_fraction__5[3], xbs_fraction__5[4], xbs_fraction__5[5], xbs_fraction__5[6], xbs_fraction__5[7], xbs_fraction__5[8], xbs_fraction__5[9], xbs_fraction__5[10], xbs_fraction__5[11], xbs_fraction__5[12], xbs_fraction__5[13], xbs_fraction__5[14], xbs_fraction__5[15], xbs_fraction__5[16], xbs_fraction__5[17], xbs_fraction__5[18], xbs_fraction__5[19], xbs_fraction__5[20], xbs_fraction__5[21], xbs_fraction__5[22], xbs_fraction__5[23], xbs_fraction__5[24], xbs_fraction__5[25], xbs_fraction__5[26], xbs_fraction__5[27]};
  assign one_hot_164291 = {reverse_164283[27:0] == 28'h000_0000, reverse_164283[27] && reverse_164283[26:0] == 27'h000_0000, reverse_164283[26] && reverse_164283[25:0] == 26'h000_0000, reverse_164283[25] && reverse_164283[24:0] == 25'h000_0000, reverse_164283[24] && reverse_164283[23:0] == 24'h00_0000, reverse_164283[23] && reverse_164283[22:0] == 23'h00_0000, reverse_164283[22] && reverse_164283[21:0] == 22'h00_0000, reverse_164283[21] && reverse_164283[20:0] == 21'h00_0000, reverse_164283[20] && reverse_164283[19:0] == 20'h0_0000, reverse_164283[19] && reverse_164283[18:0] == 19'h0_0000, reverse_164283[18] && reverse_164283[17:0] == 18'h0_0000, reverse_164283[17] && reverse_164283[16:0] == 17'h0_0000, reverse_164283[16] && reverse_164283[15:0] == 16'h0000, reverse_164283[15] && reverse_164283[14:0] == 15'h0000, reverse_164283[14] && reverse_164283[13:0] == 14'h0000, reverse_164283[13] && reverse_164283[12:0] == 13'h0000, reverse_164283[12] && reverse_164283[11:0] == 12'h000, reverse_164283[11] && reverse_164283[10:0] == 11'h000, reverse_164283[10] && reverse_164283[9:0] == 10'h000, reverse_164283[9] && reverse_164283[8:0] == 9'h000, reverse_164283[8] && reverse_164283[7:0] == 8'h00, reverse_164283[7] && reverse_164283[6:0] == 7'h00, reverse_164283[6] && reverse_164283[5:0] == 6'h00, reverse_164283[5] && reverse_164283[4:0] == 5'h00, reverse_164283[4] && reverse_164283[3:0] == 4'h0, reverse_164283[3] && reverse_164283[2:0] == 3'h0, reverse_164283[2] && reverse_164283[1:0] == 2'h0, reverse_164283[1] && !reverse_164283[0], reverse_164283[0]};
  assign reverse_164292 = {xbs_fraction__28[0], xbs_fraction__28[1], xbs_fraction__28[2], xbs_fraction__28[3], xbs_fraction__28[4], xbs_fraction__28[5], xbs_fraction__28[6], xbs_fraction__28[7], xbs_fraction__28[8], xbs_fraction__28[9], xbs_fraction__28[10], xbs_fraction__28[11], xbs_fraction__28[12], xbs_fraction__28[13], xbs_fraction__28[14], xbs_fraction__28[15], xbs_fraction__28[16], xbs_fraction__28[17], xbs_fraction__28[18], xbs_fraction__28[19], xbs_fraction__28[20], xbs_fraction__28[21], xbs_fraction__28[22], xbs_fraction__28[23], xbs_fraction__28[24], xbs_fraction__28[25], xbs_fraction__28[26], xbs_fraction__28[27]};
  assign one_hot_164293 = {reverse_164285[27:0] == 28'h000_0000, reverse_164285[27] && reverse_164285[26:0] == 27'h000_0000, reverse_164285[26] && reverse_164285[25:0] == 26'h000_0000, reverse_164285[25] && reverse_164285[24:0] == 25'h000_0000, reverse_164285[24] && reverse_164285[23:0] == 24'h00_0000, reverse_164285[23] && reverse_164285[22:0] == 23'h00_0000, reverse_164285[22] && reverse_164285[21:0] == 22'h00_0000, reverse_164285[21] && reverse_164285[20:0] == 21'h00_0000, reverse_164285[20] && reverse_164285[19:0] == 20'h0_0000, reverse_164285[19] && reverse_164285[18:0] == 19'h0_0000, reverse_164285[18] && reverse_164285[17:0] == 18'h0_0000, reverse_164285[17] && reverse_164285[16:0] == 17'h0_0000, reverse_164285[16] && reverse_164285[15:0] == 16'h0000, reverse_164285[15] && reverse_164285[14:0] == 15'h0000, reverse_164285[14] && reverse_164285[13:0] == 14'h0000, reverse_164285[13] && reverse_164285[12:0] == 13'h0000, reverse_164285[12] && reverse_164285[11:0] == 12'h000, reverse_164285[11] && reverse_164285[10:0] == 11'h000, reverse_164285[10] && reverse_164285[9:0] == 10'h000, reverse_164285[9] && reverse_164285[8:0] == 9'h000, reverse_164285[8] && reverse_164285[7:0] == 8'h00, reverse_164285[7] && reverse_164285[6:0] == 7'h00, reverse_164285[6] && reverse_164285[5:0] == 6'h00, reverse_164285[5] && reverse_164285[4:0] == 5'h00, reverse_164285[4] && reverse_164285[3:0] == 4'h0, reverse_164285[3] && reverse_164285[2:0] == 3'h0, reverse_164285[2] && reverse_164285[1:0] == 2'h0, reverse_164285[1] && !reverse_164285[0], reverse_164285[0]};
  assign reverse_164294 = {xbs_fraction__46[0], xbs_fraction__46[1], xbs_fraction__46[2], xbs_fraction__46[3], xbs_fraction__46[4], xbs_fraction__46[5], xbs_fraction__46[6], xbs_fraction__46[7], xbs_fraction__46[8], xbs_fraction__46[9], xbs_fraction__46[10], xbs_fraction__46[11], xbs_fraction__46[12], xbs_fraction__46[13], xbs_fraction__46[14], xbs_fraction__46[15], xbs_fraction__46[16], xbs_fraction__46[17], xbs_fraction__46[18], xbs_fraction__46[19], xbs_fraction__46[20], xbs_fraction__46[21], xbs_fraction__46[22], xbs_fraction__46[23], xbs_fraction__46[24], xbs_fraction__46[25], xbs_fraction__46[26], xbs_fraction__46[27]};
  assign one_hot_164295 = {reverse_164287[27:0] == 28'h000_0000, reverse_164287[27] && reverse_164287[26:0] == 27'h000_0000, reverse_164287[26] && reverse_164287[25:0] == 26'h000_0000, reverse_164287[25] && reverse_164287[24:0] == 25'h000_0000, reverse_164287[24] && reverse_164287[23:0] == 24'h00_0000, reverse_164287[23] && reverse_164287[22:0] == 23'h00_0000, reverse_164287[22] && reverse_164287[21:0] == 22'h00_0000, reverse_164287[21] && reverse_164287[20:0] == 21'h00_0000, reverse_164287[20] && reverse_164287[19:0] == 20'h0_0000, reverse_164287[19] && reverse_164287[18:0] == 19'h0_0000, reverse_164287[18] && reverse_164287[17:0] == 18'h0_0000, reverse_164287[17] && reverse_164287[16:0] == 17'h0_0000, reverse_164287[16] && reverse_164287[15:0] == 16'h0000, reverse_164287[15] && reverse_164287[14:0] == 15'h0000, reverse_164287[14] && reverse_164287[13:0] == 14'h0000, reverse_164287[13] && reverse_164287[12:0] == 13'h0000, reverse_164287[12] && reverse_164287[11:0] == 12'h000, reverse_164287[11] && reverse_164287[10:0] == 11'h000, reverse_164287[10] && reverse_164287[9:0] == 10'h000, reverse_164287[9] && reverse_164287[8:0] == 9'h000, reverse_164287[8] && reverse_164287[7:0] == 8'h00, reverse_164287[7] && reverse_164287[6:0] == 7'h00, reverse_164287[6] && reverse_164287[5:0] == 6'h00, reverse_164287[5] && reverse_164287[4:0] == 5'h00, reverse_164287[4] && reverse_164287[3:0] == 4'h0, reverse_164287[3] && reverse_164287[2:0] == 3'h0, reverse_164287[2] && reverse_164287[1:0] == 2'h0, reverse_164287[1] && !reverse_164287[0], reverse_164287[0]};
  assign reverse_164296 = {xbs_fraction__64[0], xbs_fraction__64[1], xbs_fraction__64[2], xbs_fraction__64[3], xbs_fraction__64[4], xbs_fraction__64[5], xbs_fraction__64[6], xbs_fraction__64[7], xbs_fraction__64[8], xbs_fraction__64[9], xbs_fraction__64[10], xbs_fraction__64[11], xbs_fraction__64[12], xbs_fraction__64[13], xbs_fraction__64[14], xbs_fraction__64[15], xbs_fraction__64[16], xbs_fraction__64[17], xbs_fraction__64[18], xbs_fraction__64[19], xbs_fraction__64[20], xbs_fraction__64[21], xbs_fraction__64[22], xbs_fraction__64[23], xbs_fraction__64[24], xbs_fraction__64[25], xbs_fraction__64[26], xbs_fraction__64[27]};
  assign one_hot_164297 = {reverse_164289[27:0] == 28'h000_0000, reverse_164289[27] && reverse_164289[26:0] == 27'h000_0000, reverse_164289[26] && reverse_164289[25:0] == 26'h000_0000, reverse_164289[25] && reverse_164289[24:0] == 25'h000_0000, reverse_164289[24] && reverse_164289[23:0] == 24'h00_0000, reverse_164289[23] && reverse_164289[22:0] == 23'h00_0000, reverse_164289[22] && reverse_164289[21:0] == 22'h00_0000, reverse_164289[21] && reverse_164289[20:0] == 21'h00_0000, reverse_164289[20] && reverse_164289[19:0] == 20'h0_0000, reverse_164289[19] && reverse_164289[18:0] == 19'h0_0000, reverse_164289[18] && reverse_164289[17:0] == 18'h0_0000, reverse_164289[17] && reverse_164289[16:0] == 17'h0_0000, reverse_164289[16] && reverse_164289[15:0] == 16'h0000, reverse_164289[15] && reverse_164289[14:0] == 15'h0000, reverse_164289[14] && reverse_164289[13:0] == 14'h0000, reverse_164289[13] && reverse_164289[12:0] == 13'h0000, reverse_164289[12] && reverse_164289[11:0] == 12'h000, reverse_164289[11] && reverse_164289[10:0] == 11'h000, reverse_164289[10] && reverse_164289[9:0] == 10'h000, reverse_164289[9] && reverse_164289[8:0] == 9'h000, reverse_164289[8] && reverse_164289[7:0] == 8'h00, reverse_164289[7] && reverse_164289[6:0] == 7'h00, reverse_164289[6] && reverse_164289[5:0] == 6'h00, reverse_164289[5] && reverse_164289[4:0] == 5'h00, reverse_164289[4] && reverse_164289[3:0] == 4'h0, reverse_164289[3] && reverse_164289[2:0] == 3'h0, reverse_164289[2] && reverse_164289[1:0] == 2'h0, reverse_164289[1] && !reverse_164289[0], reverse_164289[0]};
  assign one_hot_164298 = {reverse_164290[27:0] == 28'h000_0000, reverse_164290[27] && reverse_164290[26:0] == 27'h000_0000, reverse_164290[26] && reverse_164290[25:0] == 26'h000_0000, reverse_164290[25] && reverse_164290[24:0] == 25'h000_0000, reverse_164290[24] && reverse_164290[23:0] == 24'h00_0000, reverse_164290[23] && reverse_164290[22:0] == 23'h00_0000, reverse_164290[22] && reverse_164290[21:0] == 22'h00_0000, reverse_164290[21] && reverse_164290[20:0] == 21'h00_0000, reverse_164290[20] && reverse_164290[19:0] == 20'h0_0000, reverse_164290[19] && reverse_164290[18:0] == 19'h0_0000, reverse_164290[18] && reverse_164290[17:0] == 18'h0_0000, reverse_164290[17] && reverse_164290[16:0] == 17'h0_0000, reverse_164290[16] && reverse_164290[15:0] == 16'h0000, reverse_164290[15] && reverse_164290[14:0] == 15'h0000, reverse_164290[14] && reverse_164290[13:0] == 14'h0000, reverse_164290[13] && reverse_164290[12:0] == 13'h0000, reverse_164290[12] && reverse_164290[11:0] == 12'h000, reverse_164290[11] && reverse_164290[10:0] == 11'h000, reverse_164290[10] && reverse_164290[9:0] == 10'h000, reverse_164290[9] && reverse_164290[8:0] == 9'h000, reverse_164290[8] && reverse_164290[7:0] == 8'h00, reverse_164290[7] && reverse_164290[6:0] == 7'h00, reverse_164290[6] && reverse_164290[5:0] == 6'h00, reverse_164290[5] && reverse_164290[4:0] == 5'h00, reverse_164290[4] && reverse_164290[3:0] == 4'h0, reverse_164290[3] && reverse_164290[2:0] == 3'h0, reverse_164290[2] && reverse_164290[1:0] == 2'h0, reverse_164290[1] && !reverse_164290[0], reverse_164290[0]};
  assign encode_164299 = {one_hot_164291[16] | one_hot_164291[17] | one_hot_164291[18] | one_hot_164291[19] | one_hot_164291[20] | one_hot_164291[21] | one_hot_164291[22] | one_hot_164291[23] | one_hot_164291[24] | one_hot_164291[25] | one_hot_164291[26] | one_hot_164291[27] | one_hot_164291[28], one_hot_164291[8] | one_hot_164291[9] | one_hot_164291[10] | one_hot_164291[11] | one_hot_164291[12] | one_hot_164291[13] | one_hot_164291[14] | one_hot_164291[15] | one_hot_164291[24] | one_hot_164291[25] | one_hot_164291[26] | one_hot_164291[27] | one_hot_164291[28], one_hot_164291[4] | one_hot_164291[5] | one_hot_164291[6] | one_hot_164291[7] | one_hot_164291[12] | one_hot_164291[13] | one_hot_164291[14] | one_hot_164291[15] | one_hot_164291[20] | one_hot_164291[21] | one_hot_164291[22] | one_hot_164291[23] | one_hot_164291[28], one_hot_164291[2] | one_hot_164291[3] | one_hot_164291[6] | one_hot_164291[7] | one_hot_164291[10] | one_hot_164291[11] | one_hot_164291[14] | one_hot_164291[15] | one_hot_164291[18] | one_hot_164291[19] | one_hot_164291[22] | one_hot_164291[23] | one_hot_164291[26] | one_hot_164291[27], one_hot_164291[1] | one_hot_164291[3] | one_hot_164291[5] | one_hot_164291[7] | one_hot_164291[9] | one_hot_164291[11] | one_hot_164291[13] | one_hot_164291[15] | one_hot_164291[17] | one_hot_164291[19] | one_hot_164291[21] | one_hot_164291[23] | one_hot_164291[25] | one_hot_164291[27]};
  assign one_hot_164300 = {reverse_164292[27:0] == 28'h000_0000, reverse_164292[27] && reverse_164292[26:0] == 27'h000_0000, reverse_164292[26] && reverse_164292[25:0] == 26'h000_0000, reverse_164292[25] && reverse_164292[24:0] == 25'h000_0000, reverse_164292[24] && reverse_164292[23:0] == 24'h00_0000, reverse_164292[23] && reverse_164292[22:0] == 23'h00_0000, reverse_164292[22] && reverse_164292[21:0] == 22'h00_0000, reverse_164292[21] && reverse_164292[20:0] == 21'h00_0000, reverse_164292[20] && reverse_164292[19:0] == 20'h0_0000, reverse_164292[19] && reverse_164292[18:0] == 19'h0_0000, reverse_164292[18] && reverse_164292[17:0] == 18'h0_0000, reverse_164292[17] && reverse_164292[16:0] == 17'h0_0000, reverse_164292[16] && reverse_164292[15:0] == 16'h0000, reverse_164292[15] && reverse_164292[14:0] == 15'h0000, reverse_164292[14] && reverse_164292[13:0] == 14'h0000, reverse_164292[13] && reverse_164292[12:0] == 13'h0000, reverse_164292[12] && reverse_164292[11:0] == 12'h000, reverse_164292[11] && reverse_164292[10:0] == 11'h000, reverse_164292[10] && reverse_164292[9:0] == 10'h000, reverse_164292[9] && reverse_164292[8:0] == 9'h000, reverse_164292[8] && reverse_164292[7:0] == 8'h00, reverse_164292[7] && reverse_164292[6:0] == 7'h00, reverse_164292[6] && reverse_164292[5:0] == 6'h00, reverse_164292[5] && reverse_164292[4:0] == 5'h00, reverse_164292[4] && reverse_164292[3:0] == 4'h0, reverse_164292[3] && reverse_164292[2:0] == 3'h0, reverse_164292[2] && reverse_164292[1:0] == 2'h0, reverse_164292[1] && !reverse_164292[0], reverse_164292[0]};
  assign encode_164301 = {one_hot_164293[16] | one_hot_164293[17] | one_hot_164293[18] | one_hot_164293[19] | one_hot_164293[20] | one_hot_164293[21] | one_hot_164293[22] | one_hot_164293[23] | one_hot_164293[24] | one_hot_164293[25] | one_hot_164293[26] | one_hot_164293[27] | one_hot_164293[28], one_hot_164293[8] | one_hot_164293[9] | one_hot_164293[10] | one_hot_164293[11] | one_hot_164293[12] | one_hot_164293[13] | one_hot_164293[14] | one_hot_164293[15] | one_hot_164293[24] | one_hot_164293[25] | one_hot_164293[26] | one_hot_164293[27] | one_hot_164293[28], one_hot_164293[4] | one_hot_164293[5] | one_hot_164293[6] | one_hot_164293[7] | one_hot_164293[12] | one_hot_164293[13] | one_hot_164293[14] | one_hot_164293[15] | one_hot_164293[20] | one_hot_164293[21] | one_hot_164293[22] | one_hot_164293[23] | one_hot_164293[28], one_hot_164293[2] | one_hot_164293[3] | one_hot_164293[6] | one_hot_164293[7] | one_hot_164293[10] | one_hot_164293[11] | one_hot_164293[14] | one_hot_164293[15] | one_hot_164293[18] | one_hot_164293[19] | one_hot_164293[22] | one_hot_164293[23] | one_hot_164293[26] | one_hot_164293[27], one_hot_164293[1] | one_hot_164293[3] | one_hot_164293[5] | one_hot_164293[7] | one_hot_164293[9] | one_hot_164293[11] | one_hot_164293[13] | one_hot_164293[15] | one_hot_164293[17] | one_hot_164293[19] | one_hot_164293[21] | one_hot_164293[23] | one_hot_164293[25] | one_hot_164293[27]};
  assign one_hot_164302 = {reverse_164294[27:0] == 28'h000_0000, reverse_164294[27] && reverse_164294[26:0] == 27'h000_0000, reverse_164294[26] && reverse_164294[25:0] == 26'h000_0000, reverse_164294[25] && reverse_164294[24:0] == 25'h000_0000, reverse_164294[24] && reverse_164294[23:0] == 24'h00_0000, reverse_164294[23] && reverse_164294[22:0] == 23'h00_0000, reverse_164294[22] && reverse_164294[21:0] == 22'h00_0000, reverse_164294[21] && reverse_164294[20:0] == 21'h00_0000, reverse_164294[20] && reverse_164294[19:0] == 20'h0_0000, reverse_164294[19] && reverse_164294[18:0] == 19'h0_0000, reverse_164294[18] && reverse_164294[17:0] == 18'h0_0000, reverse_164294[17] && reverse_164294[16:0] == 17'h0_0000, reverse_164294[16] && reverse_164294[15:0] == 16'h0000, reverse_164294[15] && reverse_164294[14:0] == 15'h0000, reverse_164294[14] && reverse_164294[13:0] == 14'h0000, reverse_164294[13] && reverse_164294[12:0] == 13'h0000, reverse_164294[12] && reverse_164294[11:0] == 12'h000, reverse_164294[11] && reverse_164294[10:0] == 11'h000, reverse_164294[10] && reverse_164294[9:0] == 10'h000, reverse_164294[9] && reverse_164294[8:0] == 9'h000, reverse_164294[8] && reverse_164294[7:0] == 8'h00, reverse_164294[7] && reverse_164294[6:0] == 7'h00, reverse_164294[6] && reverse_164294[5:0] == 6'h00, reverse_164294[5] && reverse_164294[4:0] == 5'h00, reverse_164294[4] && reverse_164294[3:0] == 4'h0, reverse_164294[3] && reverse_164294[2:0] == 3'h0, reverse_164294[2] && reverse_164294[1:0] == 2'h0, reverse_164294[1] && !reverse_164294[0], reverse_164294[0]};
  assign encode_164303 = {one_hot_164295[16] | one_hot_164295[17] | one_hot_164295[18] | one_hot_164295[19] | one_hot_164295[20] | one_hot_164295[21] | one_hot_164295[22] | one_hot_164295[23] | one_hot_164295[24] | one_hot_164295[25] | one_hot_164295[26] | one_hot_164295[27] | one_hot_164295[28], one_hot_164295[8] | one_hot_164295[9] | one_hot_164295[10] | one_hot_164295[11] | one_hot_164295[12] | one_hot_164295[13] | one_hot_164295[14] | one_hot_164295[15] | one_hot_164295[24] | one_hot_164295[25] | one_hot_164295[26] | one_hot_164295[27] | one_hot_164295[28], one_hot_164295[4] | one_hot_164295[5] | one_hot_164295[6] | one_hot_164295[7] | one_hot_164295[12] | one_hot_164295[13] | one_hot_164295[14] | one_hot_164295[15] | one_hot_164295[20] | one_hot_164295[21] | one_hot_164295[22] | one_hot_164295[23] | one_hot_164295[28], one_hot_164295[2] | one_hot_164295[3] | one_hot_164295[6] | one_hot_164295[7] | one_hot_164295[10] | one_hot_164295[11] | one_hot_164295[14] | one_hot_164295[15] | one_hot_164295[18] | one_hot_164295[19] | one_hot_164295[22] | one_hot_164295[23] | one_hot_164295[26] | one_hot_164295[27], one_hot_164295[1] | one_hot_164295[3] | one_hot_164295[5] | one_hot_164295[7] | one_hot_164295[9] | one_hot_164295[11] | one_hot_164295[13] | one_hot_164295[15] | one_hot_164295[17] | one_hot_164295[19] | one_hot_164295[21] | one_hot_164295[23] | one_hot_164295[25] | one_hot_164295[27]};
  assign one_hot_164304 = {reverse_164296[27:0] == 28'h000_0000, reverse_164296[27] && reverse_164296[26:0] == 27'h000_0000, reverse_164296[26] && reverse_164296[25:0] == 26'h000_0000, reverse_164296[25] && reverse_164296[24:0] == 25'h000_0000, reverse_164296[24] && reverse_164296[23:0] == 24'h00_0000, reverse_164296[23] && reverse_164296[22:0] == 23'h00_0000, reverse_164296[22] && reverse_164296[21:0] == 22'h00_0000, reverse_164296[21] && reverse_164296[20:0] == 21'h00_0000, reverse_164296[20] && reverse_164296[19:0] == 20'h0_0000, reverse_164296[19] && reverse_164296[18:0] == 19'h0_0000, reverse_164296[18] && reverse_164296[17:0] == 18'h0_0000, reverse_164296[17] && reverse_164296[16:0] == 17'h0_0000, reverse_164296[16] && reverse_164296[15:0] == 16'h0000, reverse_164296[15] && reverse_164296[14:0] == 15'h0000, reverse_164296[14] && reverse_164296[13:0] == 14'h0000, reverse_164296[13] && reverse_164296[12:0] == 13'h0000, reverse_164296[12] && reverse_164296[11:0] == 12'h000, reverse_164296[11] && reverse_164296[10:0] == 11'h000, reverse_164296[10] && reverse_164296[9:0] == 10'h000, reverse_164296[9] && reverse_164296[8:0] == 9'h000, reverse_164296[8] && reverse_164296[7:0] == 8'h00, reverse_164296[7] && reverse_164296[6:0] == 7'h00, reverse_164296[6] && reverse_164296[5:0] == 6'h00, reverse_164296[5] && reverse_164296[4:0] == 5'h00, reverse_164296[4] && reverse_164296[3:0] == 4'h0, reverse_164296[3] && reverse_164296[2:0] == 3'h0, reverse_164296[2] && reverse_164296[1:0] == 2'h0, reverse_164296[1] && !reverse_164296[0], reverse_164296[0]};
  assign encode_164305 = {one_hot_164297[16] | one_hot_164297[17] | one_hot_164297[18] | one_hot_164297[19] | one_hot_164297[20] | one_hot_164297[21] | one_hot_164297[22] | one_hot_164297[23] | one_hot_164297[24] | one_hot_164297[25] | one_hot_164297[26] | one_hot_164297[27] | one_hot_164297[28], one_hot_164297[8] | one_hot_164297[9] | one_hot_164297[10] | one_hot_164297[11] | one_hot_164297[12] | one_hot_164297[13] | one_hot_164297[14] | one_hot_164297[15] | one_hot_164297[24] | one_hot_164297[25] | one_hot_164297[26] | one_hot_164297[27] | one_hot_164297[28], one_hot_164297[4] | one_hot_164297[5] | one_hot_164297[6] | one_hot_164297[7] | one_hot_164297[12] | one_hot_164297[13] | one_hot_164297[14] | one_hot_164297[15] | one_hot_164297[20] | one_hot_164297[21] | one_hot_164297[22] | one_hot_164297[23] | one_hot_164297[28], one_hot_164297[2] | one_hot_164297[3] | one_hot_164297[6] | one_hot_164297[7] | one_hot_164297[10] | one_hot_164297[11] | one_hot_164297[14] | one_hot_164297[15] | one_hot_164297[18] | one_hot_164297[19] | one_hot_164297[22] | one_hot_164297[23] | one_hot_164297[26] | one_hot_164297[27], one_hot_164297[1] | one_hot_164297[3] | one_hot_164297[5] | one_hot_164297[7] | one_hot_164297[9] | one_hot_164297[11] | one_hot_164297[13] | one_hot_164297[15] | one_hot_164297[17] | one_hot_164297[19] | one_hot_164297[21] | one_hot_164297[23] | one_hot_164297[25] | one_hot_164297[27]};
  assign encode_164306 = {one_hot_164298[16] | one_hot_164298[17] | one_hot_164298[18] | one_hot_164298[19] | one_hot_164298[20] | one_hot_164298[21] | one_hot_164298[22] | one_hot_164298[23] | one_hot_164298[24] | one_hot_164298[25] | one_hot_164298[26] | one_hot_164298[27] | one_hot_164298[28], one_hot_164298[8] | one_hot_164298[9] | one_hot_164298[10] | one_hot_164298[11] | one_hot_164298[12] | one_hot_164298[13] | one_hot_164298[14] | one_hot_164298[15] | one_hot_164298[24] | one_hot_164298[25] | one_hot_164298[26] | one_hot_164298[27] | one_hot_164298[28], one_hot_164298[4] | one_hot_164298[5] | one_hot_164298[6] | one_hot_164298[7] | one_hot_164298[12] | one_hot_164298[13] | one_hot_164298[14] | one_hot_164298[15] | one_hot_164298[20] | one_hot_164298[21] | one_hot_164298[22] | one_hot_164298[23] | one_hot_164298[28], one_hot_164298[2] | one_hot_164298[3] | one_hot_164298[6] | one_hot_164298[7] | one_hot_164298[10] | one_hot_164298[11] | one_hot_164298[14] | one_hot_164298[15] | one_hot_164298[18] | one_hot_164298[19] | one_hot_164298[22] | one_hot_164298[23] | one_hot_164298[26] | one_hot_164298[27], one_hot_164298[1] | one_hot_164298[3] | one_hot_164298[5] | one_hot_164298[7] | one_hot_164298[9] | one_hot_164298[11] | one_hot_164298[13] | one_hot_164298[15] | one_hot_164298[17] | one_hot_164298[19] | one_hot_164298[21] | one_hot_164298[23] | one_hot_164298[25] | one_hot_164298[27]};
  assign encode_164308 = {one_hot_164300[16] | one_hot_164300[17] | one_hot_164300[18] | one_hot_164300[19] | one_hot_164300[20] | one_hot_164300[21] | one_hot_164300[22] | one_hot_164300[23] | one_hot_164300[24] | one_hot_164300[25] | one_hot_164300[26] | one_hot_164300[27] | one_hot_164300[28], one_hot_164300[8] | one_hot_164300[9] | one_hot_164300[10] | one_hot_164300[11] | one_hot_164300[12] | one_hot_164300[13] | one_hot_164300[14] | one_hot_164300[15] | one_hot_164300[24] | one_hot_164300[25] | one_hot_164300[26] | one_hot_164300[27] | one_hot_164300[28], one_hot_164300[4] | one_hot_164300[5] | one_hot_164300[6] | one_hot_164300[7] | one_hot_164300[12] | one_hot_164300[13] | one_hot_164300[14] | one_hot_164300[15] | one_hot_164300[20] | one_hot_164300[21] | one_hot_164300[22] | one_hot_164300[23] | one_hot_164300[28], one_hot_164300[2] | one_hot_164300[3] | one_hot_164300[6] | one_hot_164300[7] | one_hot_164300[10] | one_hot_164300[11] | one_hot_164300[14] | one_hot_164300[15] | one_hot_164300[18] | one_hot_164300[19] | one_hot_164300[22] | one_hot_164300[23] | one_hot_164300[26] | one_hot_164300[27], one_hot_164300[1] | one_hot_164300[3] | one_hot_164300[5] | one_hot_164300[7] | one_hot_164300[9] | one_hot_164300[11] | one_hot_164300[13] | one_hot_164300[15] | one_hot_164300[17] | one_hot_164300[19] | one_hot_164300[21] | one_hot_164300[23] | one_hot_164300[25] | one_hot_164300[27]};
  assign encode_164310 = {one_hot_164302[16] | one_hot_164302[17] | one_hot_164302[18] | one_hot_164302[19] | one_hot_164302[20] | one_hot_164302[21] | one_hot_164302[22] | one_hot_164302[23] | one_hot_164302[24] | one_hot_164302[25] | one_hot_164302[26] | one_hot_164302[27] | one_hot_164302[28], one_hot_164302[8] | one_hot_164302[9] | one_hot_164302[10] | one_hot_164302[11] | one_hot_164302[12] | one_hot_164302[13] | one_hot_164302[14] | one_hot_164302[15] | one_hot_164302[24] | one_hot_164302[25] | one_hot_164302[26] | one_hot_164302[27] | one_hot_164302[28], one_hot_164302[4] | one_hot_164302[5] | one_hot_164302[6] | one_hot_164302[7] | one_hot_164302[12] | one_hot_164302[13] | one_hot_164302[14] | one_hot_164302[15] | one_hot_164302[20] | one_hot_164302[21] | one_hot_164302[22] | one_hot_164302[23] | one_hot_164302[28], one_hot_164302[2] | one_hot_164302[3] | one_hot_164302[6] | one_hot_164302[7] | one_hot_164302[10] | one_hot_164302[11] | one_hot_164302[14] | one_hot_164302[15] | one_hot_164302[18] | one_hot_164302[19] | one_hot_164302[22] | one_hot_164302[23] | one_hot_164302[26] | one_hot_164302[27], one_hot_164302[1] | one_hot_164302[3] | one_hot_164302[5] | one_hot_164302[7] | one_hot_164302[9] | one_hot_164302[11] | one_hot_164302[13] | one_hot_164302[15] | one_hot_164302[17] | one_hot_164302[19] | one_hot_164302[21] | one_hot_164302[23] | one_hot_164302[25] | one_hot_164302[27]};
  assign encode_164312 = {one_hot_164304[16] | one_hot_164304[17] | one_hot_164304[18] | one_hot_164304[19] | one_hot_164304[20] | one_hot_164304[21] | one_hot_164304[22] | one_hot_164304[23] | one_hot_164304[24] | one_hot_164304[25] | one_hot_164304[26] | one_hot_164304[27] | one_hot_164304[28], one_hot_164304[8] | one_hot_164304[9] | one_hot_164304[10] | one_hot_164304[11] | one_hot_164304[12] | one_hot_164304[13] | one_hot_164304[14] | one_hot_164304[15] | one_hot_164304[24] | one_hot_164304[25] | one_hot_164304[26] | one_hot_164304[27] | one_hot_164304[28], one_hot_164304[4] | one_hot_164304[5] | one_hot_164304[6] | one_hot_164304[7] | one_hot_164304[12] | one_hot_164304[13] | one_hot_164304[14] | one_hot_164304[15] | one_hot_164304[20] | one_hot_164304[21] | one_hot_164304[22] | one_hot_164304[23] | one_hot_164304[28], one_hot_164304[2] | one_hot_164304[3] | one_hot_164304[6] | one_hot_164304[7] | one_hot_164304[10] | one_hot_164304[11] | one_hot_164304[14] | one_hot_164304[15] | one_hot_164304[18] | one_hot_164304[19] | one_hot_164304[22] | one_hot_164304[23] | one_hot_164304[26] | one_hot_164304[27], one_hot_164304[1] | one_hot_164304[3] | one_hot_164304[5] | one_hot_164304[7] | one_hot_164304[9] | one_hot_164304[11] | one_hot_164304[13] | one_hot_164304[15] | one_hot_164304[17] | one_hot_164304[19] | one_hot_164304[21] | one_hot_164304[23] | one_hot_164304[25] | one_hot_164304[27]};
  assign cancel__14 = |encode_164299[4:1];
  assign carry_bit__13 = xbs_fraction__13[27];
  assign result_fraction__502 = 23'h00_0000;
  assign cancel__28 = |encode_164301[4:1];
  assign carry_bit__28 = xbs_fraction__27[27];
  assign result_fraction__569 = 23'h00_0000;
  assign cancel__47 = |encode_164303[4:1];
  assign carry_bit__47 = xbs_fraction__45[27];
  assign result_fraction__634 = 23'h00_0000;
  assign cancel__66 = |encode_164305[4:1];
  assign carry_bit__66 = xbs_fraction__63[27];
  assign result_fraction__707 = 23'h00_0000;
  assign cancel__5 = |encode_164306[4:1];
  assign carry_bit__5 = xbs_fraction__5[27];
  assign result_fraction__503 = 23'h00_0000;
  assign leading_zeroes__13 = {result_fraction__502, encode_164299};
  assign cancel__29 = |encode_164308[4:1];
  assign carry_bit__29 = xbs_fraction__28[27];
  assign result_fraction__570 = 23'h00_0000;
  assign leading_zeroes__28 = {result_fraction__569, encode_164301};
  assign cancel__48 = |encode_164310[4:1];
  assign carry_bit__48 = xbs_fraction__46[27];
  assign result_fraction__635 = 23'h00_0000;
  assign leading_zeroes__47 = {result_fraction__634, encode_164303};
  assign cancel__67 = |encode_164312[4:1];
  assign carry_bit__67 = xbs_fraction__64[27];
  assign result_fraction__708 = 23'h00_0000;
  assign leading_zeroes__66 = {result_fraction__707, encode_164305};
  assign leading_zeroes__5 = {result_fraction__503, encode_164306};
  assign carry_fraction__26 = xbs_fraction__13[27:1];
  assign add_164379 = leading_zeroes__13 + 28'hfff_ffff;
  assign leading_zeroes__29 = {result_fraction__570, encode_164308};
  assign carry_fraction__55 = xbs_fraction__27[27:1];
  assign add_164392 = leading_zeroes__28 + 28'hfff_ffff;
  assign leading_zeroes__48 = {result_fraction__635, encode_164310};
  assign carry_fraction__93 = xbs_fraction__45[27:1];
  assign add_164405 = leading_zeroes__47 + 28'hfff_ffff;
  assign leading_zeroes__67 = {result_fraction__708, encode_164312};
  assign array_index_164412 = in_img_unflattened[4'hb];
  assign carry_fraction__131 = xbs_fraction__63[27:1];
  assign add_164419 = leading_zeroes__66 + 28'hfff_ffff;
  assign carry_fraction__9 = xbs_fraction__5[27:1];
  assign add_164426 = leading_zeroes__5 + 28'hfff_ffff;
  assign concat_164427 = {~(carry_bit__13 | cancel__14), ~(carry_bit__13 | ~cancel__14), ~(~carry_bit__13 | cancel__14)};
  assign carry_fraction__27 = carry_fraction__26 | {26'h000_0000, xbs_fraction__13[0]};
  assign cancel_fraction__13 = add_164379 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__13[26:0] << add_164379;
  assign carry_fraction__56 = xbs_fraction__28[27:1];
  assign add_164436 = leading_zeroes__29 + 28'hfff_ffff;
  assign concat_164437 = {~(carry_bit__28 | cancel__28), ~(carry_bit__28 | ~cancel__28), ~(~carry_bit__28 | cancel__28)};
  assign carry_fraction__57 = carry_fraction__55 | {26'h000_0000, xbs_fraction__27[0]};
  assign cancel_fraction__28 = add_164392 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__27[26:0] << add_164392;
  assign carry_fraction__94 = xbs_fraction__46[27:1];
  assign add_164446 = leading_zeroes__48 + 28'hfff_ffff;
  assign concat_164447 = {~(carry_bit__47 | cancel__47), ~(carry_bit__47 | ~cancel__47), ~(~carry_bit__47 | cancel__47)};
  assign carry_fraction__95 = carry_fraction__93 | {26'h000_0000, xbs_fraction__45[0]};
  assign cancel_fraction__47 = add_164405 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__45[26:0] << add_164405;
  assign carry_fraction__132 = xbs_fraction__64[27:1];
  assign add_164456 = leading_zeroes__67 + 28'hfff_ffff;
  assign x_bexp__510 = array_index_164412[30:23];
  assign concat_164458 = {~(carry_bit__66 | cancel__66), ~(carry_bit__66 | ~cancel__66), ~(~carry_bit__66 | cancel__66)};
  assign carry_fraction__133 = carry_fraction__131 | {26'h000_0000, xbs_fraction__63[0]};
  assign cancel_fraction__66 = add_164419 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__63[26:0] << add_164419;
  assign concat_164461 = {~(carry_bit__5 | cancel__5), ~(carry_bit__5 | ~cancel__5), ~(~carry_bit__5 | cancel__5)};
  assign carry_fraction__10 = carry_fraction__9 | {26'h000_0000, xbs_fraction__5[0]};
  assign cancel_fraction__5 = add_164426 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__5[26:0] << add_164426;
  assign shifted_fraction__13 = carry_fraction__27 & {27{concat_164427[0]}} | cancel_fraction__13 & {27{concat_164427[1]}} | xbs_fraction__13[26:0] & {27{concat_164427[2]}};
  assign concat_164465 = {~(carry_bit__29 | cancel__29), ~(carry_bit__29 | ~cancel__29), ~(~carry_bit__29 | cancel__29)};
  assign carry_fraction__58 = carry_fraction__56 | {26'h000_0000, xbs_fraction__28[0]};
  assign cancel_fraction__29 = add_164436 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__28[26:0] << add_164436;
  assign result_sign__1023 = 1'h0;
  assign shifted_fraction__28 = carry_fraction__57 & {27{concat_164437[0]}} | cancel_fraction__28 & {27{concat_164437[1]}} | xbs_fraction__27[26:0] & {27{concat_164437[2]}};
  assign concat_164471 = {~(carry_bit__48 | cancel__48), ~(carry_bit__48 | ~cancel__48), ~(~carry_bit__48 | cancel__48)};
  assign carry_fraction__96 = carry_fraction__94 | {26'h000_0000, xbs_fraction__46[0]};
  assign cancel_fraction__48 = add_164446 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__46[26:0] << add_164446;
  assign result_sign__1024 = 1'h0;
  assign shifted_fraction__47 = carry_fraction__95 & {27{concat_164447[0]}} | cancel_fraction__47 & {27{concat_164447[1]}} | xbs_fraction__45[26:0] & {27{concat_164447[2]}};
  assign concat_164477 = {~(carry_bit__67 | cancel__67), ~(carry_bit__67 | ~cancel__67), ~(~carry_bit__67 | cancel__67)};
  assign carry_fraction__134 = carry_fraction__132 | {26'h000_0000, xbs_fraction__64[0]};
  assign cancel_fraction__67 = add_164456 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__64[26:0] << add_164456;
  assign result_sign__1025 = 1'h0;
  assign shifted_fraction__66 = carry_fraction__133 & {27{concat_164458[0]}} | cancel_fraction__66 & {27{concat_164458[1]}} | xbs_fraction__63[26:0] & {27{concat_164458[2]}};
  assign shifted_fraction__5 = carry_fraction__10 & {27{concat_164461[0]}} | cancel_fraction__5 & {27{concat_164461[1]}} | xbs_fraction__5[26:0] & {27{concat_164461[2]}};
  assign result_sign__1026 = 1'h0;
  assign shifted_fraction__29 = carry_fraction__58 & {27{concat_164465[0]}} | cancel_fraction__29 & {27{concat_164465[1]}} | xbs_fraction__28[26:0] & {27{concat_164465[2]}};
  assign result_sign__1027 = 1'h0;
  assign shifted_fraction__48 = carry_fraction__96 & {27{concat_164471[0]}} | cancel_fraction__48 & {27{concat_164471[1]}} | xbs_fraction__46[26:0] & {27{concat_164471[2]}};
  assign result_sign__1028 = 1'h0;
  assign shifted_fraction__67 = carry_fraction__134 & {27{concat_164477[0]}} | cancel_fraction__67 & {27{concat_164477[1]}} | xbs_fraction__64[26:0] & {27{concat_164477[2]}};
  assign result_sign__1029 = 1'h0;
  assign result_sign__1030 = 1'h0;
  assign normal_chunk__13 = shifted_fraction__13[2:0];
  assign fraction_shift__241 = 3'h4;
  assign half_way_chunk__13 = shifted_fraction__13[3:2];
  assign result_sign__1031 = 1'h0;
  assign result_sign__1107 = 1'h0;
  assign add_164512 = {result_sign__1023, x_bexp__461[7]} + 2'h1;
  assign normal_chunk__28 = shifted_fraction__28[2:0];
  assign fraction_shift__276 = 3'h4;
  assign half_way_chunk__28 = shifted_fraction__28[3:2];
  assign result_sign__1032 = 1'h0;
  assign result_sign__1110 = 1'h0;
  assign add_164523 = {result_sign__1024, x_bexp__503[7]} + 2'h1;
  assign x_bexp__742 = 8'h00;
  assign result_sign__616 = 1'h0;
  assign x_fraction__505 = array_index_163484[22:0];
  assign normal_chunk__47 = shifted_fraction__47[2:0];
  assign fraction_shift__311 = 3'h4;
  assign half_way_chunk__47 = shifted_fraction__47[3:2];
  assign result_sign__1033 = 1'h0;
  assign result_sign__1114 = 1'h0;
  assign add_164537 = {result_sign__1025, x_bexp__510[7]} + 2'h1;
  assign x_bexp__743 = 8'h00;
  assign result_sign__723 = 1'h0;
  assign x_fraction__510 = array_index_164412[22:0];
  assign normal_chunk__66 = shifted_fraction__66[2:0];
  assign fraction_shift__346 = 3'h4;
  assign half_way_chunk__66 = shifted_fraction__66[3:2];
  assign normal_chunk__5 = shifted_fraction__5[2:0];
  assign fraction_shift__242 = 3'h4;
  assign half_way_chunk__5 = shifted_fraction__5[3:2];
  assign result_sign__424 = 1'h0;
  assign add_164557 = {result_sign__1026, shifted_fraction__13[26:3]} + 25'h000_0001;
  assign normal_chunk__29 = shifted_fraction__29[2:0];
  assign fraction_shift__277 = 3'h4;
  assign half_way_chunk__29 = shifted_fraction__29[3:2];
  assign result_sign__519 = 1'h0;
  assign add_164569 = {result_sign__1027, shifted_fraction__28[26:3]} + 25'h000_0001;
  assign normal_chunk__48 = shifted_fraction__48[2:0];
  assign fraction_shift__312 = 3'h4;
  assign half_way_chunk__48 = shifted_fraction__48[3:2];
  assign ne_164578 = x_bexp__503 != x_bexp__742;
  assign result_sign__618 = 1'h0;
  assign add_164584 = {result_sign__1028, shifted_fraction__47[26:3]} + 25'h000_0001;
  assign normal_chunk__67 = shifted_fraction__67[2:0];
  assign fraction_shift__347 = 3'h4;
  assign half_way_chunk__67 = shifted_fraction__67[3:2];
  assign ne_164593 = x_bexp__510 != x_bexp__743;
  assign result_sign__725 = 1'h0;
  assign add_164599 = {result_sign__1029, shifted_fraction__66[26:3]} + 25'h000_0001;
  assign result_sign__425 = 1'h0;
  assign add_164603 = {result_sign__1030, shifted_fraction__5[26:3]} + 25'h000_0001;
  assign do_round_up__27 = normal_chunk__13 > fraction_shift__241 | half_way_chunk__13 == 2'h3;
  assign result_sign__520 = 1'h0;
  assign add_164610 = {result_sign__1031, shifted_fraction__29[26:3]} + 25'h000_0001;
  assign exp__124 = {result_sign__1107, add_164512, x_bexp__461[6:0]} + 10'h381;
  assign do_round_up__58 = normal_chunk__28 > fraction_shift__276 | half_way_chunk__28 == 2'h3;
  assign result_sign__619 = 1'h0;
  assign add_164618 = {result_sign__1032, shifted_fraction__48[26:3]} + 25'h000_0001;
  assign exp__206 = {result_sign__1110, add_164523, x_bexp__503[6:0]} + 10'h381;
  assign sign_ext_164620 = {10{ne_164578}};
  assign x_fraction__368 = {result_sign__616, x_fraction__505} | 24'h80_0000;
  assign do_round_up__97 = normal_chunk__47 > fraction_shift__311 | half_way_chunk__47 == 2'h3;
  assign result_sign__726 = 1'h0;
  assign add_164629 = {result_sign__1033, shifted_fraction__67[26:3]} + 25'h000_0001;
  assign exp__288 = {result_sign__1114, add_164537, x_bexp__510[6:0]} + 10'h381;
  assign sign_ext_164631 = {10{ne_164593}};
  assign x_fraction__512 = {result_sign__723, x_fraction__510} | 24'h80_0000;
  assign do_round_up__136 = normal_chunk__66 > fraction_shift__346 | half_way_chunk__66 == 2'h3;
  assign do_round_up__10 = normal_chunk__5 > fraction_shift__242 | half_way_chunk__5 == 2'h3;
  assign rounded_fraction__13 = do_round_up__27 ? {add_164557, normal_chunk__13} : {result_sign__424, shifted_fraction__13};
  assign do_round_up__59 = normal_chunk__29 > fraction_shift__277 | half_way_chunk__29 == 2'h3;
  assign exp__126 = exp__124 & sign_ext_159707;
  assign rounded_fraction__28 = do_round_up__58 ? {add_164569, normal_chunk__28} : {result_sign__519, shifted_fraction__28};
  assign do_round_up__98 = normal_chunk__48 > fraction_shift__312 | half_way_chunk__48 == 2'h3;
  assign exp__208 = exp__206 & sign_ext_164620;
  assign x_fraction__370 = x_fraction__368 & {24{ne_164578}};
  assign result_sign__816 = 1'h0;
  assign result_sign__817 = 1'h0;
  assign rounded_fraction__47 = do_round_up__97 ? {add_164584, normal_chunk__47} : {result_sign__618, shifted_fraction__47};
  assign do_round_up__137 = normal_chunk__67 > fraction_shift__347 | half_way_chunk__67 == 2'h3;
  assign exp__290 = exp__288 & sign_ext_164631;
  assign x_fraction__514 = x_fraction__512 & {24{ne_164593}};
  assign result_sign__818 = 1'h0;
  assign result_sign__819 = 1'h0;
  assign rounded_fraction__66 = do_round_up__136 ? {add_164599, normal_chunk__66} : {result_sign__725, shifted_fraction__66};
  assign rounded_fraction__5 = do_round_up__10 ? {add_164603, normal_chunk__5} : {result_sign__425, shifted_fraction__5};
  assign result_sign__426 = 1'h0;
  assign x_bexp__582 = 8'h00;
  assign rounding_carry__13 = rounded_fraction__13[27];
  assign rounded_fraction__29 = do_round_up__59 ? {add_164610, normal_chunk__29} : {result_sign__520, shifted_fraction__29};
  assign result_sign__521 = 1'h0;
  assign x_bexp__600 = 8'h00;
  assign rounding_carry__28 = rounded_fraction__28[27];
  assign rounded_fraction__48 = do_round_up__98 ? {add_164618, normal_chunk__48} : {result_sign__619, shifted_fraction__48};
  assign concat_164676 = {x_fraction__370, result_sign__816};
  assign concat_164677 = {result_sign__817, x_fraction__370};
  assign result_sign__620 = 1'h0;
  assign x_bexp__618 = 8'h00;
  assign rounding_carry__47 = rounded_fraction__47[27];
  assign rounded_fraction__67 = do_round_up__137 ? {add_164629, normal_chunk__67} : {result_sign__726, shifted_fraction__67};
  assign concat_164683 = {x_fraction__514, result_sign__818};
  assign concat_164684 = {result_sign__819, x_fraction__514};
  assign result_sign__727 = 1'h0;
  assign x_bexp__636 = 8'h00;
  assign rounding_carry__66 = rounded_fraction__66[27];
  assign result_sign__427 = 1'h0;
  assign x_bexp__583 = 8'h00;
  assign rounding_carry__5 = rounded_fraction__5[27];
  assign result_sign__522 = 1'h0;
  assign x_bexp__601 = 8'h00;
  assign rounding_carry__29 = rounded_fraction__29[27];
  assign sel_164696 = $signed(exp__126) <= $signed(10'h000) ? concat_159775 : concat_159774;
  assign result_sign__621 = 1'h0;
  assign x_bexp__619 = 8'h00;
  assign rounding_carry__48 = rounded_fraction__48[27];
  assign sel_164702 = $signed(exp__208) <= $signed(10'h000) ? concat_164677 : concat_164676;
  assign result_sign__728 = 1'h0;
  assign x_bexp__637 = 8'h00;
  assign rounding_carry__67 = rounded_fraction__67[27];
  assign sel_164708 = $signed(exp__290) <= $signed(10'h000) ? concat_164684 : concat_164683;
  assign result_sign__428 = 1'h0;
  assign add_164714 = {result_sign__426, x_bexp__110} + {x_bexp__582, rounding_carry__13};
  assign result_sign__937 = 1'h0;
  assign fraction__281 = sel_164696[23:1];
  assign result_sign__523 = 1'h0;
  assign add_164722 = {result_sign__521, x_bexp__219} + {x_bexp__600, rounding_carry__28};
  assign result_sign__944 = 1'h0;
  assign fraction__460 = sel_164702[23:1];
  assign result_sign__622 = 1'h0;
  assign add_164730 = {result_sign__620, x_bexp__363} + {x_bexp__618, rounding_carry__47};
  assign result_sign__952 = 1'h0;
  assign fraction__639 = sel_164708[23:1];
  assign result_sign__729 = 1'h0;
  assign add_164738 = {result_sign__727, x_bexp__507} + {x_bexp__636, rounding_carry__66};
  assign result_sign__429 = 1'h0;
  assign add_164742 = {result_sign__427, x_bexp__38} + {x_bexp__583, rounding_carry__5};
  assign result_sign__524 = 1'h0;
  assign add_164751 = {result_sign__522, x_bexp__220} + {x_bexp__601, rounding_carry__29};
  assign fraction__283 = {result_sign__937, fraction__281};
  assign result_sign__623 = 1'h0;
  assign add_164764 = {result_sign__621, x_bexp__364} + {x_bexp__619, rounding_carry__48};
  assign fraction__462 = {result_sign__944, fraction__460};
  assign result_sign__730 = 1'h0;
  assign add_164777 = {result_sign__728, x_bexp__508} + {x_bexp__637, rounding_carry__67};
  assign fraction__641 = {result_sign__952, fraction__639};
  assign add_164794 = {result_sign__428, add_164714} + 10'h001;
  assign do_round_up__61 = sel_164696[0] & sel_164696[1];
  assign add_164803 = fraction__283 + 24'h00_0001;
  assign add_164804 = {result_sign__523, add_164722} + 10'h001;
  assign do_round_up__100 = sel_164702[0] & sel_164702[1];
  assign add_164813 = fraction__462 + 24'h00_0001;
  assign add_164814 = {result_sign__622, add_164730} + 10'h001;
  assign do_round_up__139 = sel_164708[0] & sel_164708[1];
  assign add_164823 = fraction__641 + 24'h00_0001;
  assign add_164824 = {result_sign__729, add_164738} + 10'h001;
  assign add_164827 = {result_sign__429, add_164742} + 10'h001;
  assign wide_exponent__39 = add_164794 - {5'h00, encode_164299};
  assign add_164832 = {result_sign__524, add_164751} + 10'h001;
  assign fraction__285 = do_round_up__61 ? add_164803 : fraction__283;
  assign wide_exponent__82 = add_164804 - {5'h00, encode_164301};
  assign add_164839 = {result_sign__623, add_164764} + 10'h001;
  assign fraction__464 = do_round_up__100 ? add_164813 : fraction__462;
  assign wide_exponent__139 = add_164814 - {5'h00, encode_164303};
  assign add_164846 = {result_sign__730, add_164777} + 10'h001;
  assign fraction__643 = do_round_up__139 ? add_164823 : fraction__641;
  assign wide_exponent__196 = add_164824 - {5'h00, encode_164305};
  assign wide_exponent__13 = add_164827 - {5'h00, encode_164306};
  assign wide_exponent__40 = wide_exponent__39 & {10{add_164224 != 26'h000_0000 | xddend_y__13[2:0] != 3'h0}};
  assign wide_exponent__83 = add_164832 - {5'h00, encode_164308};
  assign add_164859 = exp__126 + 10'h001;
  assign wide_exponent__84 = wide_exponent__82 & {10{add_164227 != 26'h000_0000 | xddend_y__27[2:0] != 3'h0}};
  assign wide_exponent__140 = add_164839 - {5'h00, encode_164310};
  assign add_164864 = exp__208 + 10'h001;
  assign wide_exponent__141 = wide_exponent__139 & {10{add_164230 != 26'h000_0000 | xddend_y__45[2:0] != 3'h0}};
  assign wide_exponent__197 = add_164846 - {5'h00, encode_164312};
  assign add_164869 = exp__290 + 10'h001;
  assign wide_exponent__198 = wide_exponent__196 & {10{add_164233 != 26'h000_0000 | xddend_y__63[2:0] != 3'h0}};
  assign wide_exponent__14 = wide_exponent__13 & {10{add_164234 != 26'h000_0000 | xddend_y__5[2:0] != 3'h0}};
  assign high_exp__371 = 8'hff;
  assign result_fraction__777 = 23'h00_0000;
  assign high_exp__372 = 8'hff;
  assign result_fraction__778 = 23'h00_0000;
  assign high_exp__104 = 8'hff;
  assign result_fraction__504 = 23'h00_0000;
  assign high_exp__105 = 8'hff;
  assign result_fraction__505 = 23'h00_0000;
  assign wide_exponent__85 = wide_exponent__83 & {10{add_164237 != 26'h000_0000 | xddend_y__28[2:0] != 3'h0}};
  assign exp__130 = fraction__285[23] ? add_164859 : exp__126;
  assign high_exp__403 = 8'hff;
  assign result_fraction__810 = 23'h00_0000;
  assign high_exp__404 = 8'hff;
  assign result_fraction__811 = 23'h00_0000;
  assign high_exp__168 = 8'hff;
  assign result_fraction__571 = 23'h00_0000;
  assign high_exp__169 = 8'hff;
  assign result_fraction__572 = 23'h00_0000;
  assign wide_exponent__142 = wide_exponent__140 & {10{add_164240 != 26'h000_0000 | xddend_y__46[2:0] != 3'h0}};
  assign exp__212 = fraction__464[23] ? add_164864 : exp__208;
  assign high_exp__435 = 8'hff;
  assign result_fraction__843 = 23'h00_0000;
  assign high_exp__436 = 8'hff;
  assign result_fraction__844 = 23'h00_0000;
  assign high_exp__234 = 8'hff;
  assign result_fraction__636 = 23'h00_0000;
  assign high_exp__235 = 8'hff;
  assign result_fraction__637 = 23'h00_0000;
  assign wide_exponent__199 = wide_exponent__197 & {10{add_164243 != 26'h000_0000 | xddend_y__64[2:0] != 3'h0}};
  assign exp__294 = fraction__643[23] ? add_164869 : exp__290;
  assign high_exp__467 = 8'hff;
  assign result_fraction__876 = 23'h00_0000;
  assign high_exp__468 = 8'hff;
  assign result_fraction__877 = 23'h00_0000;
  assign high_exp__305 = 8'hff;
  assign result_fraction__709 = 23'h00_0000;
  assign high_exp__306 = 8'hff;
  assign result_fraction__710 = 23'h00_0000;
  assign high_exp__357 = 8'hff;
  assign result_fraction__762 = 23'h00_0000;
  assign high_exp__358 = 8'hff;
  assign result_fraction__763 = 23'h00_0000;
  assign high_exp__106 = 8'hff;
  assign result_fraction__506 = 23'h00_0000;
  assign high_exp__107 = 8'hff;
  assign result_fraction__507 = 23'h00_0000;
  assign ne_164928 = x_fraction__110 != result_fraction__777;
  assign ne_164930 = prod_fraction__39 != result_fraction__778;
  assign eq_164931 = x_bexp__110 == high_exp__104;
  assign eq_164932 = x_fraction__110 == result_fraction__504;
  assign eq_164933 = prod_bexp__54 == high_exp__105;
  assign eq_164934 = prod_fraction__39 == result_fraction__505;
  assign high_exp__389 = 8'hff;
  assign result_fraction__795 = 23'h00_0000;
  assign high_exp__390 = 8'hff;
  assign result_fraction__796 = 23'h00_0000;
  assign high_exp__170 = 8'hff;
  assign result_fraction__573 = 23'h00_0000;
  assign high_exp__171 = 8'hff;
  assign result_fraction__574 = 23'h00_0000;
  assign ne_164947 = x_fraction__219 != result_fraction__810;
  assign ne_164949 = prod_fraction__79 != result_fraction__811;
  assign eq_164950 = x_bexp__219 == high_exp__168;
  assign eq_164951 = x_fraction__219 == result_fraction__571;
  assign eq_164952 = prod_bexp__107 == high_exp__169;
  assign eq_164953 = prod_fraction__79 == result_fraction__572;
  assign high_exp__421 = 8'hff;
  assign result_fraction__828 = 23'h00_0000;
  assign high_exp__422 = 8'hff;
  assign result_fraction__829 = 23'h00_0000;
  assign high_exp__236 = 8'hff;
  assign result_fraction__638 = 23'h00_0000;
  assign high_exp__237 = 8'hff;
  assign result_fraction__639 = 23'h00_0000;
  assign ne_164966 = x_fraction__363 != result_fraction__843;
  assign ne_164968 = prod_fraction__133 != result_fraction__844;
  assign eq_164969 = x_bexp__363 == high_exp__234;
  assign eq_164970 = x_fraction__363 == result_fraction__636;
  assign eq_164971 = prod_bexp__179 == high_exp__235;
  assign eq_164972 = prod_fraction__133 == result_fraction__637;
  assign high_exp__453 = 8'hff;
  assign result_fraction__861 = 23'h00_0000;
  assign high_exp__454 = 8'hff;
  assign result_fraction__862 = 23'h00_0000;
  assign high_exp__307 = 8'hff;
  assign result_fraction__711 = 23'h00_0000;
  assign high_exp__308 = 8'hff;
  assign result_fraction__712 = 23'h00_0000;
  assign ne_164985 = x_fraction__507 != result_fraction__876;
  assign ne_164987 = prod_fraction__187 != result_fraction__877;
  assign eq_164988 = x_bexp__507 == high_exp__305;
  assign eq_164989 = x_fraction__507 == result_fraction__709;
  assign eq_164990 = prod_bexp__251 == high_exp__306;
  assign eq_164991 = prod_fraction__187 == result_fraction__710;
  assign ne_164994 = x_fraction__38 != result_fraction__762;
  assign ne_164996 = prod_fraction__13 != result_fraction__763;
  assign eq_164997 = x_bexp__38 == high_exp__106;
  assign eq_164998 = x_fraction__38 == result_fraction__506;
  assign eq_164999 = prod_bexp__18 == high_exp__107;
  assign eq_165000 = prod_fraction__13 == result_fraction__507;
  assign ne_165009 = x_fraction__220 != result_fraction__795;
  assign ne_165011 = prod_fraction__80 != result_fraction__796;
  assign eq_165012 = x_bexp__220 == high_exp__170;
  assign eq_165013 = x_fraction__220 == result_fraction__573;
  assign eq_165014 = prod_bexp__108 == high_exp__171;
  assign eq_165015 = prod_fraction__80 == result_fraction__574;
  assign result_exp__92 = exp__130[8:0];
  assign ne_165026 = x_fraction__364 != result_fraction__828;
  assign ne_165028 = prod_fraction__134 != result_fraction__829;
  assign eq_165029 = x_bexp__364 == high_exp__236;
  assign eq_165030 = x_fraction__364 == result_fraction__638;
  assign eq_165031 = prod_bexp__180 == high_exp__237;
  assign eq_165032 = prod_fraction__134 == result_fraction__639;
  assign result_exp__152 = exp__212[8:0];
  assign ne_165043 = x_fraction__508 != result_fraction__861;
  assign ne_165045 = prod_fraction__188 != result_fraction__862;
  assign eq_165046 = x_bexp__508 == high_exp__307;
  assign eq_165047 = x_fraction__508 == result_fraction__711;
  assign eq_165048 = prod_bexp__252 == high_exp__308;
  assign eq_165049 = prod_fraction__188 == result_fraction__712;
  assign result_exp__212 = exp__294[8:0];
  assign wide_exponent__41 = wide_exponent__40[8:0] & {9{~wide_exponent__40[9]}};
  assign has_pos_inf__13 = ~(x_bexp__110 != high_exp__371 | ne_164928 | x_sign__28) | ~(prod_bexp__54 != high_exp__372 | ne_164930 | prod_sign__13);
  assign has_neg_inf__13 = eq_164931 & eq_164932 & x_sign__28 | eq_164933 & eq_164934 & prod_sign__13;
  assign result_exp__94 = result_exp__92 & {9{$signed(exp__130) > $signed(10'h000)}};
  assign wide_exponent__86 = wide_exponent__84[8:0] & {9{~wide_exponent__84[9]}};
  assign has_pos_inf__28 = ~(x_bexp__219 != high_exp__403 | ne_164947 | x_sign__55) | ~(prod_bexp__107 != high_exp__404 | ne_164949 | prod_sign__27);
  assign has_neg_inf__28 = eq_164950 & eq_164951 & x_sign__55 | eq_164952 & eq_164953 & prod_sign__27;
  assign result_fraction__706 = 23'h00_0000;
  assign result_fraction__705 = 23'h00_0000;
  assign result_exp__154 = result_exp__152 & {9{$signed(exp__212) > $signed(10'h000)}};
  assign wide_exponent__143 = wide_exponent__141[8:0] & {9{~wide_exponent__141[9]}};
  assign has_pos_inf__47 = ~(x_bexp__363 != high_exp__435 | ne_164966 | x_sign__91) | ~(prod_bexp__179 != high_exp__436 | ne_164968 | prod_sign__45);
  assign has_neg_inf__47 = eq_164969 & eq_164970 & x_sign__91 | eq_164971 & eq_164972 & prod_sign__45;
  assign high_exp__310 = 8'hff;
  assign result_fraction__714 = 23'h00_0000;
  assign result_fraction__713 = 23'h00_0000;
  assign result_exp__214 = result_exp__212 & {9{$signed(exp__294) > $signed(10'h000)}};
  assign wide_exponent__200 = wide_exponent__198[8:0] & {9{~wide_exponent__198[9]}};
  assign has_pos_inf__66 = ~(x_bexp__507 != high_exp__467 | ne_164985 | x_sign__127) | ~(prod_bexp__251 != high_exp__468 | ne_164987 | prod_sign__63);
  assign has_neg_inf__66 = eq_164988 & eq_164989 & x_sign__127 | eq_164990 & eq_164991 & prod_sign__63;
  assign wide_exponent__15 = wide_exponent__14[8:0] & {9{~wide_exponent__14[9]}};
  assign has_pos_inf__5 = ~(x_bexp__38 != high_exp__357 | ne_164994 | x_sign__10) | ~(prod_bexp__18 != high_exp__358 | ne_164996 | prod_sign__5);
  assign has_neg_inf__5 = eq_164997 & eq_164998 & x_sign__10 | eq_164999 & eq_165000 & prod_sign__5;
  assign wide_exponent__87 = wide_exponent__85[8:0] & {9{~wide_exponent__85[9]}};
  assign has_pos_inf__29 = ~(x_bexp__220 != high_exp__389 | ne_165009 | x_sign__56) | ~(prod_bexp__108 != high_exp__390 | ne_165011 | prod_sign__28);
  assign has_neg_inf__29 = eq_165012 & eq_165013 & x_sign__56 | eq_165014 & eq_165015 & prod_sign__28;
  assign wide_exponent__144 = wide_exponent__142[8:0] & {9{~wide_exponent__142[9]}};
  assign has_pos_inf__48 = ~(x_bexp__364 != high_exp__421 | ne_165026 | x_sign__92) | ~(prod_bexp__180 != high_exp__422 | ne_165028 | prod_sign__46);
  assign has_neg_inf__48 = eq_165029 & eq_165030 & x_sign__92 | eq_165031 & eq_165032 & prod_sign__46;
  assign ne_165126 = x_fraction__505 != result_fraction__706;
  assign wide_exponent__201 = wide_exponent__199[8:0] & {9{~wide_exponent__199[9]}};
  assign has_pos_inf__67 = ~(x_bexp__508 != high_exp__453 | ne_165043 | x_sign__128) | ~(prod_bexp__252 != high_exp__454 | ne_165045 | prod_sign__64);
  assign has_neg_inf__67 = eq_165046 & eq_165047 & x_sign__128 | eq_165048 & eq_165049 & prod_sign__64;
  assign is_result_nan__138 = x_bexp__510 == high_exp__310;
  assign ne_165140 = x_fraction__510 != result_fraction__714;
  assign is_result_nan__27 = eq_164931 & ne_164928 | eq_164933 & ne_164930 | has_pos_inf__13 & has_neg_inf__13;
  assign is_operand_inf__13 = eq_164931 & eq_164932 | eq_164933 & eq_164934;
  assign and_reduce_165162 = &wide_exponent__41[7:0];
  assign and_reduce_165171 = &result_exp__94[7:0];
  assign is_result_nan__58 = eq_164950 & ne_164947 | eq_164952 & ne_164949 | has_pos_inf__28 & has_neg_inf__28;
  assign is_operand_inf__28 = eq_164950 & eq_164951 | eq_164952 & eq_164953;
  assign and_reduce_165177 = &wide_exponent__86[7:0];
  assign is_result_nan__100 = is_result_nan__134 & ne_165126;
  assign has_inf_arg__69 = is_result_nan__134 & x_fraction__505 == result_fraction__705;
  assign and_reduce_165188 = &result_exp__154[7:0];
  assign is_result_nan__97 = eq_164969 & ne_164966 | eq_164971 & ne_164968 | has_pos_inf__47 & has_neg_inf__47;
  assign is_operand_inf__47 = eq_164969 & eq_164970 | eq_164971 & eq_164972;
  assign and_reduce_165194 = &wide_exponent__143[7:0];
  assign is_result_nan__139 = is_result_nan__138 & ne_165140;
  assign has_inf_arg__71 = is_result_nan__138 & x_fraction__510 == result_fraction__713;
  assign and_reduce_165205 = &result_exp__214[7:0];
  assign is_result_nan__136 = eq_164988 & ne_164985 | eq_164990 & ne_164987 | has_pos_inf__66 & has_neg_inf__66;
  assign is_operand_inf__66 = eq_164988 & eq_164989 | eq_164990 & eq_164991;
  assign and_reduce_165211 = &wide_exponent__200[7:0];
  assign is_result_nan__10 = eq_164997 & ne_164994 | eq_164999 & ne_164996 | has_pos_inf__5 & has_neg_inf__5;
  assign is_operand_inf__5 = eq_164997 & eq_164998 | eq_164999 & eq_165000;
  assign and_reduce_165217 = &wide_exponent__15[7:0];
  assign fraction_shift__374 = 3'h3;
  assign fraction_shift__243 = 3'h4;
  assign high_exp__108 = 8'hff;
  assign is_result_nan__59 = eq_165012 & ne_165009 | eq_165014 & ne_165011 | has_pos_inf__29 & has_neg_inf__29;
  assign is_operand_inf__29 = eq_165012 & eq_165013 | eq_165014 & eq_165015;
  assign and_reduce_165229 = &wide_exponent__87[7:0];
  assign high_exp__174 = 8'hff;
  assign fraction_shift__392 = 3'h3;
  assign fraction_shift__278 = 3'h4;
  assign high_exp__172 = 8'hff;
  assign result_exp__95 = {8{is_result_nan__60}};
  assign is_result_nan__98 = eq_165029 & ne_165026 | eq_165031 & ne_165028 | has_pos_inf__48 & has_neg_inf__48;
  assign is_operand_inf__48 = eq_165029 & eq_165030 | eq_165031 & eq_165032;
  assign and_reduce_165244 = &wide_exponent__144[7:0];
  assign high_exp__240 = 8'hff;
  assign fraction_shift__410 = 3'h3;
  assign fraction_shift__313 = 3'h4;
  assign high_exp__238 = 8'hff;
  assign is_result_nan__137 = eq_165046 & ne_165043 | eq_165048 & ne_165045 | has_pos_inf__67 & has_neg_inf__67;
  assign is_operand_inf__67 = eq_165046 & eq_165047 | eq_165048 & eq_165049;
  assign and_reduce_165258 = &wide_exponent__201[7:0];
  assign high_exp__312 = 8'hff;
  assign fraction_shift__428 = 3'h3;
  assign fraction_shift__348 = 3'h4;
  assign high_exp__309 = 8'hff;
  assign result_exp__215 = {8{is_result_nan__138}};
  assign fraction_shift__375 = 3'h3;
  assign fraction_shift__244 = 3'h4;
  assign high_exp__109 = 8'hff;
  assign fraction_shift__42 = rounding_carry__13 ? fraction_shift__243 : fraction_shift__374;
  assign result_sign__430 = 1'h0;
  assign result_exponent__14 = is_result_nan__27 | is_operand_inf__13 | wide_exponent__41[8] | and_reduce_165162 ? high_exp__108 : wide_exponent__41[7:0];
  assign fraction_shift__393 = 3'h3;
  assign fraction_shift__279 = 3'h4;
  assign is_subnormal__32 = $signed(exp__130) <= $signed(10'h000);
  assign high_exp__173 = 8'hff;
  assign result_exp__96 = is_result_nan__126 | has_inf_arg__65 | result_exp__94[8] | and_reduce_165171 ? high_exp__174 : result_exp__94[7:0];
  assign fraction_shift__86 = rounding_carry__28 ? fraction_shift__278 : fraction_shift__392;
  assign result_sign__525 = 1'h0;
  assign result_exponent__28 = is_result_nan__58 | is_operand_inf__28 | wide_exponent__86[8] | and_reduce_165177 ? high_exp__172 : wide_exponent__86[7:0];
  assign result_sign__526 = 1'h0;
  assign fraction_shift__411 = 3'h3;
  assign fraction_shift__314 = 3'h4;
  assign is_subnormal__52 = $signed(exp__212) <= $signed(10'h000);
  assign high_exp__239 = 8'hff;
  assign result_exp__156 = is_result_nan__100 | has_inf_arg__69 | result_exp__154[8] | and_reduce_165188 ? high_exp__240 : result_exp__154[7:0];
  assign fraction_shift__143 = rounding_carry__47 ? fraction_shift__313 : fraction_shift__410;
  assign result_sign__624 = 1'h0;
  assign result_exponent__47 = is_result_nan__97 | is_operand_inf__47 | wide_exponent__143[8] | and_reduce_165194 ? high_exp__238 : wide_exponent__143[7:0];
  assign fraction_shift__429 = 3'h3;
  assign fraction_shift__349 = 3'h4;
  assign is_subnormal__72 = $signed(exp__294) <= $signed(10'h000);
  assign high_exp__311 = 8'hff;
  assign result_exp__216 = is_result_nan__139 | has_inf_arg__71 | result_exp__214[8] | and_reduce_165205 ? high_exp__312 : result_exp__214[7:0];
  assign fraction_shift__200 = rounding_carry__66 ? fraction_shift__348 : fraction_shift__428;
  assign result_sign__731 = 1'h0;
  assign result_exponent__66 = is_result_nan__136 | is_operand_inf__66 | wide_exponent__200[8] | and_reduce_165211 ? high_exp__309 : wide_exponent__200[7:0];
  assign result_sign__732 = 1'h0;
  assign fraction_shift__15 = rounding_carry__5 ? fraction_shift__244 : fraction_shift__375;
  assign result_sign__431 = 1'h0;
  assign result_exponent__5 = is_result_nan__10 | is_operand_inf__5 | wide_exponent__15[8] | and_reduce_165217 ? high_exp__109 : wide_exponent__15[7:0];
  assign shrl_165317 = rounded_fraction__13 >> fraction_shift__42;
  assign fraction_shift__87 = rounding_carry__29 ? fraction_shift__279 : fraction_shift__393;
  assign result_sign__527 = 1'h0;
  assign result_exponent__29 = is_result_nan__59 | is_operand_inf__29 | wide_exponent__87[8] | and_reduce_165229 ? high_exp__173 : wide_exponent__87[7:0];
  assign result_sign__528 = 1'h0;
  assign shrl_165327 = rounded_fraction__28 >> fraction_shift__86;
  assign fraction_shift__144 = rounding_carry__48 ? fraction_shift__314 : fraction_shift__411;
  assign result_sign__625 = 1'h0;
  assign result_exponent__48 = is_result_nan__98 | is_operand_inf__48 | wide_exponent__144[8] | and_reduce_165244 ? high_exp__239 : wide_exponent__144[7:0];
  assign result_sign__626 = 1'h0;
  assign shrl_165338 = rounded_fraction__47 >> fraction_shift__143;
  assign fraction_shift__201 = rounding_carry__67 ? fraction_shift__349 : fraction_shift__429;
  assign result_sign__733 = 1'h0;
  assign result_exponent__67 = is_result_nan__137 | is_operand_inf__67 | wide_exponent__201[8] | and_reduce_165258 ? high_exp__311 : wide_exponent__201[7:0];
  assign result_sign__734 = 1'h0;
  assign shrl_165348 = rounded_fraction__66 >> fraction_shift__200;
  assign shrl_165352 = rounded_fraction__5 >> fraction_shift__15;
  assign result_fraction__81 = shrl_165317[22:0];
  assign sum__14 = {result_sign__430, result_exponent__14} + concat_158884;
  assign shrl_165358 = rounded_fraction__29 >> fraction_shift__87;
  assign result_fraction__172 = shrl_165327[22:0];
  assign sum__30 = {result_sign__525, result_exponent__28} + {result_sign__526, ~result_exp__95};
  assign shrl_165366 = rounded_fraction__48 >> fraction_shift__144;
  assign concat_165370 = {result_sign__626, ~result_exp__156};
  assign result_fraction__289 = shrl_165338[22:0];
  assign sum__49 = {result_sign__624, result_exponent__47} + concat_163691;
  assign shrl_165374 = rounded_fraction__67 >> fraction_shift__201;
  assign result_fraction__406 = shrl_165348[22:0];
  assign sum__68 = {result_sign__731, result_exponent__66} + {result_sign__732, ~result_exp__215};
  assign result_fraction__28 = shrl_165352[22:0];
  assign sum__6 = {result_sign__431, result_exponent__5} + concat_158865;
  assign result_fraction__82 = result_fraction__81 & {23{~(is_operand_inf__13 | wide_exponent__41[8] | and_reduce_165162 | ~((|wide_exponent__41[8:1]) | wide_exponent__41[0]))}};
  assign nan_fraction__91 = 23'h40_0000;
  assign result_fraction__173 = shrl_165358[22:0];
  assign result_fraction__179 = fraction__285[22:0];
  assign sum__31 = {result_sign__527, result_exponent__29} + {result_sign__528, ~result_exp__96};
  assign result_fraction__174 = result_fraction__172 & {23{~(is_operand_inf__28 | wide_exponent__86[8] | and_reduce_165177 | ~((|wide_exponent__86[8:1]) | wide_exponent__86[0]))}};
  assign nan_fraction__117 = 23'h40_0000;
  assign result_fraction__290 = shrl_165366[22:0];
  assign result_fraction__296 = fraction__464[22:0];
  assign sum__50 = {result_sign__625, result_exponent__48} + concat_165370;
  assign result_fraction__291 = result_fraction__289 & {23{~(is_operand_inf__47 | wide_exponent__143[8] | and_reduce_165194 | ~((|wide_exponent__143[8:1]) | wide_exponent__143[0]))}};
  assign nan_fraction__145 = 23'h40_0000;
  assign result_fraction__407 = shrl_165374[22:0];
  assign result_fraction__413 = fraction__643[22:0];
  assign sum__69 = {result_sign__733, result_exponent__67} + {result_sign__734, ~result_exp__216};
  assign result_fraction__408 = result_fraction__406 & {23{~(is_operand_inf__66 | wide_exponent__200[8] | and_reduce_165211 | ~((|wide_exponent__200[8:1]) | wide_exponent__200[0]))}};
  assign nan_fraction__174 = 23'h40_0000;
  assign result_fraction__29 = result_fraction__28 & {23{~(is_operand_inf__5 | wide_exponent__15[8] | and_reduce_165217 | ~((|wide_exponent__15[8:1]) | wide_exponent__15[0]))}};
  assign nan_fraction__92 = 23'h40_0000;
  assign result_fraction__83 = is_result_nan__27 ? nan_fraction__91 : result_fraction__82;
  assign prod_bexp__58 = sum__14[8] ? result_exp__192 : result_exponent__14;
  assign x_bexp__744 = 8'h00;
  assign result_fraction__175 = result_fraction__173 & {23{~(is_operand_inf__29 | wide_exponent__87[8] | and_reduce_165229 | ~((|wide_exponent__87[8:1]) | wide_exponent__87[0]))}};
  assign nan_fraction__118 = 23'h40_0000;
  assign result_fraction__181 = result_fraction__179 & {23{~(has_inf_arg__65 | result_exp__94[8] | and_reduce_165171 | is_subnormal__32)}};
  assign nan_fraction__119 = 23'h40_0000;
  assign result_fraction__176 = is_result_nan__58 ? nan_fraction__117 : result_fraction__174;
  assign result_fraction__477 = {is_result_nan__60, 22'h00_0000};
  assign prod_bexp__115 = sum__30[8] ? result_exp__95 : result_exponent__28;
  assign x_bexp__745 = 8'h00;
  assign result_fraction__292 = result_fraction__290 & {23{~(is_operand_inf__48 | wide_exponent__144[8] | and_reduce_165244 | ~((|wide_exponent__144[8:1]) | wide_exponent__144[0]))}};
  assign nan_fraction__146 = 23'h40_0000;
  assign result_fraction__298 = result_fraction__296 & {23{~(has_inf_arg__69 | result_exp__154[8] | and_reduce_165188 | is_subnormal__52)}};
  assign nan_fraction__147 = 23'h40_0000;
  assign result_fraction__293 = is_result_nan__97 ? nan_fraction__145 : result_fraction__291;
  assign prod_bexp__187 = sum__49[8] ? result_exp__209 : result_exponent__47;
  assign x_bexp__746 = 8'h00;
  assign result_fraction__409 = result_fraction__407 & {23{~(is_operand_inf__67 | wide_exponent__201[8] | and_reduce_165258 | ~((|wide_exponent__201[8:1]) | wide_exponent__201[0]))}};
  assign nan_fraction__175 = 23'h40_0000;
  assign result_fraction__415 = result_fraction__413 & {23{~(has_inf_arg__71 | result_exp__214[8] | and_reduce_165205 | is_subnormal__72)}};
  assign nan_fraction__176 = 23'h40_0000;
  assign result_fraction__410 = is_result_nan__136 ? nan_fraction__174 : result_fraction__408;
  assign result_fraction__478 = {is_result_nan__138, 22'h00_0000};
  assign prod_bexp__259 = sum__68[8] ? result_exp__215 : result_exponent__66;
  assign x_bexp__747 = 8'h00;
  assign result_fraction__30 = is_result_nan__10 ? nan_fraction__92 : result_fraction__29;
  assign prod_bexp__22 = sum__6[8] ? result_exp__191 : result_exponent__5;
  assign x_bexp__748 = 8'h00;
  assign fraction_is_zero__13 = add_164224 == 26'h000_0000 & xddend_y__13[2:0] == 3'h0;
  assign prod_fraction__42 = sum__14[8] ? result_fraction__472 : result_fraction__83;
  assign incremented_sum__86 = sum__14[7:0] + 8'h01;
  assign result_fraction__177 = is_result_nan__59 ? nan_fraction__118 : result_fraction__175;
  assign result_fraction__183 = is_result_nan__126 ? nan_fraction__119 : result_fraction__181;
  assign prod_bexp__116 = sum__31[8] ? result_exp__96 : result_exponent__29;
  assign x_bexp__749 = 8'h00;
  assign fraction_is_zero__28 = add_164227 == 26'h000_0000 & xddend_y__27[2:0] == 3'h0;
  assign prod_fraction__85 = sum__30[8] ? result_fraction__477 : result_fraction__176;
  assign incremented_sum__104 = sum__30[7:0] + 8'h01;
  assign result_fraction__294 = is_result_nan__98 ? nan_fraction__146 : result_fraction__292;
  assign result_fraction__300 = is_result_nan__100 ? nan_fraction__147 : result_fraction__298;
  assign prod_bexp__188 = sum__50[8] ? result_exp__156 : result_exponent__48;
  assign x_bexp__750 = 8'h00;
  assign fraction_is_zero__47 = add_164230 == 26'h000_0000 & xddend_y__45[2:0] == 3'h0;
  assign prod_fraction__139 = sum__49[8] ? result_fraction__476 : result_fraction__293;
  assign incremented_sum__122 = sum__49[7:0] + 8'h01;
  assign result_fraction__411 = is_result_nan__137 ? nan_fraction__175 : result_fraction__409;
  assign result_fraction__417 = is_result_nan__139 ? nan_fraction__176 : result_fraction__415;
  assign prod_bexp__260 = sum__69[8] ? result_exp__216 : result_exponent__67;
  assign x_bexp__751 = 8'h00;
  assign fraction_is_zero__66 = add_164233 == 26'h000_0000 & xddend_y__63[2:0] == 3'h0;
  assign prod_fraction__193 = sum__68[8] ? result_fraction__478 : result_fraction__410;
  assign incremented_sum__140 = sum__68[7:0] + 8'h01;
  assign fraction_is_zero__5 = add_164234 == 26'h000_0000 & xddend_y__5[2:0] == 3'h0;
  assign prod_fraction__16 = sum__6[8] ? result_fraction__368 : result_fraction__30;
  assign incremented_sum__87 = sum__6[7:0] + 8'h01;
  assign wide_y__28 = {2'h1, prod_fraction__42, 3'h0};
  assign x_bexpbs_difference__15 = sum__14[8] ? incremented_sum__86 : ~sum__14[7:0];
  assign fraction_is_zero__29 = add_164237 == 26'h000_0000 & xddend_y__28[2:0] == 3'h0;
  assign prod_fraction__86 = sum__31[8] ? result_fraction__183 : result_fraction__177;
  assign incremented_sum__105 = sum__31[7:0] + 8'h01;
  assign wide_y__59 = {2'h1, prod_fraction__85, 3'h0};
  assign x_bexpbs_difference__29 = sum__30[8] ? incremented_sum__104 : ~sum__30[7:0];
  assign fraction_is_zero__48 = add_164240 == 26'h000_0000 & xddend_y__46[2:0] == 3'h0;
  assign prod_fraction__140 = sum__50[8] ? result_fraction__300 : result_fraction__294;
  assign incremented_sum__123 = sum__50[7:0] + 8'h01;
  assign wide_y__97 = {2'h1, prod_fraction__139, 3'h0};
  assign x_bexpbs_difference__47 = sum__49[8] ? incremented_sum__122 : ~sum__49[7:0];
  assign fraction_is_zero__67 = add_164243 == 26'h000_0000 & xddend_y__64[2:0] == 3'h0;
  assign prod_fraction__194 = sum__69[8] ? result_fraction__417 : result_fraction__411;
  assign incremented_sum__141 = sum__69[7:0] + 8'h01;
  assign wide_y__135 = {2'h1, prod_fraction__193, 3'h0};
  assign x_bexpbs_difference__65 = sum__68[8] ? incremented_sum__140 : ~sum__68[7:0];
  assign wide_y__11 = {2'h1, prod_fraction__16, 3'h0};
  assign x_bexpbs_difference__6 = sum__6[8] ? incremented_sum__87 : ~sum__6[7:0];
  assign concat_165590 = {~(add_164224[25] | fraction_is_zero__13), add_164224[25], fraction_is_zero__13};
  assign x_bexp__118 = sum__14[8] ? result_exponent__14 : result_exp__192;
  assign x_bexp__752 = 8'h00;
  assign wide_y__29 = wide_y__28 & {28{prod_bexp__58 != x_bexp__744}};
  assign sub_165596 = 8'h1c - x_bexpbs_difference__15;
  assign wide_y__60 = {2'h1, prod_fraction__86, 3'h0};
  assign x_bexpbs_difference__30 = sum__31[8] ? incremented_sum__105 : ~sum__31[7:0];
  assign concat_165602 = {~(add_164227[25] | fraction_is_zero__28), add_164227[25], fraction_is_zero__28};
  assign x_bexp__235 = sum__30[8] ? result_exponent__28 : result_exp__95;
  assign x_bexp__753 = 8'h00;
  assign wide_y__61 = wide_y__59 & {28{prod_bexp__115 != x_bexp__745}};
  assign sub_165608 = 8'h1c - x_bexpbs_difference__29;
  assign wide_y__98 = {2'h1, prod_fraction__140, 3'h0};
  assign x_bexpbs_difference__48 = sum__50[8] ? incremented_sum__123 : ~sum__50[7:0];
  assign concat_165614 = {~(add_164230[25] | fraction_is_zero__47), add_164230[25], fraction_is_zero__47};
  assign x_bexp__379 = sum__49[8] ? result_exponent__47 : result_exp__209;
  assign x_bexp__754 = 8'h00;
  assign wide_y__99 = wide_y__97 & {28{prod_bexp__187 != x_bexp__746}};
  assign sub_165620 = 8'h1c - x_bexpbs_difference__47;
  assign wide_y__136 = {2'h1, prod_fraction__194, 3'h0};
  assign x_bexpbs_difference__66 = sum__69[8] ? incremented_sum__141 : ~sum__69[7:0];
  assign concat_165626 = {~(add_164233[25] | fraction_is_zero__66), add_164233[25], fraction_is_zero__66};
  assign x_bexp__523 = sum__68[8] ? result_exponent__66 : result_exp__215;
  assign x_bexp__755 = 8'h00;
  assign wide_y__137 = wide_y__135 & {28{prod_bexp__259 != x_bexp__747}};
  assign sub_165632 = 8'h1c - x_bexpbs_difference__65;
  assign concat_165633 = {~(add_164234[25] | fraction_is_zero__5), add_164234[25], fraction_is_zero__5};
  assign x_bexp__46 = sum__6[8] ? result_exponent__5 : result_exp__191;
  assign x_bexp__756 = 8'h00;
  assign wide_y__12 = wide_y__11 & {28{prod_bexp__22 != x_bexp__748}};
  assign sub_165639 = 8'h1c - x_bexpbs_difference__6;
  assign result_sign__67 = x_sign__28 & prod_sign__13 & concat_165590[0] | ~prod_sign__13 & concat_165590[1] | prod_sign__13 & concat_165590[2];
  assign x_fraction__118 = sum__14[8] ? result_fraction__83 : result_fraction__472;
  assign dropped__14 = sub_165596 >= 8'h1c ? 28'h000_0000 : wide_y__29 << sub_165596;
  assign concat_165647 = {~(add_164237[25] | fraction_is_zero__29), add_164237[25], fraction_is_zero__29};
  assign x_bexp__236 = sum__31[8] ? result_exponent__29 : result_exp__96;
  assign x_bexp__757 = 8'h00;
  assign wide_y__62 = wide_y__60 & {28{prod_bexp__116 != x_bexp__749}};
  assign sub_165653 = 8'h1c - x_bexpbs_difference__30;
  assign high_exp__482 = 8'hff;
  assign result_sign__142 = x_sign__55 & prod_sign__27 & concat_165602[0] | ~prod_sign__27 & concat_165602[1] | prod_sign__27 & concat_165602[2];
  assign x_fraction__235 = sum__30[8] ? result_fraction__176 : result_fraction__477;
  assign dropped__30 = sub_165608 >= 8'h1c ? 28'h000_0000 : wide_y__61 << sub_165608;
  assign concat_165662 = {~(add_164240[25] | fraction_is_zero__48), add_164240[25], fraction_is_zero__48};
  assign x_bexp__380 = sum__50[8] ? result_exponent__48 : result_exp__156;
  assign x_bexp__758 = 8'h00;
  assign wide_y__100 = wide_y__98 & {28{prod_bexp__188 != x_bexp__750}};
  assign sub_165668 = 8'h1c - x_bexpbs_difference__48;
  assign result_sign__239 = x_sign__91 & prod_sign__45 & concat_165614[0] | ~prod_sign__45 & concat_165614[1] | prod_sign__45 & concat_165614[2];
  assign x_fraction__379 = sum__49[8] ? result_fraction__293 : result_fraction__476;
  assign dropped__49 = sub_165620 >= 8'h1c ? 28'h000_0000 : wide_y__99 << sub_165620;
  assign concat_165676 = {~(add_164243[25] | fraction_is_zero__67), add_164243[25], fraction_is_zero__67};
  assign x_bexp__524 = sum__69[8] ? result_exponent__67 : result_exp__216;
  assign x_bexp__759 = 8'h00;
  assign wide_y__138 = wide_y__136 & {28{prod_bexp__260 != x_bexp__751}};
  assign sub_165682 = 8'h1c - x_bexpbs_difference__66;
  assign high_exp__489 = 8'hff;
  assign result_sign__336 = x_sign__127 & prod_sign__63 & concat_165626[0] | ~prod_sign__63 & concat_165626[1] | prod_sign__63 & concat_165626[2];
  assign x_fraction__523 = sum__68[8] ? result_fraction__410 : result_fraction__478;
  assign dropped__68 = sub_165632 >= 8'h1c ? 28'h000_0000 : wide_y__137 << sub_165632;
  assign result_sign__23 = x_sign__10 & prod_sign__5 & concat_165633[0] | ~prod_sign__5 & concat_165633[1] | prod_sign__5 & concat_165633[2];
  assign x_fraction__46 = sum__6[8] ? result_fraction__30 : result_fraction__368;
  assign dropped__6 = sub_165639 >= 8'h1c ? 28'h000_0000 : wide_y__12 << sub_165639;
  assign result_sign__68 = is_operand_inf__13 ? ~has_pos_inf__13 : result_sign__67;
  assign wide_x__28 = {2'h1, x_fraction__118, 3'h0};
  assign result_sign__143 = x_sign__56 & prod_sign__28 & concat_165647[0] | ~prod_sign__28 & concat_165647[1] | prod_sign__28 & concat_165647[2];
  assign x_fraction__236 = sum__31[8] ? result_fraction__177 : result_fraction__183;
  assign dropped__31 = sub_165653 >= 8'h1c ? 28'h000_0000 : wide_y__62 << sub_165653;
  assign result_sign__144 = is_operand_inf__28 ? ~has_pos_inf__28 : result_sign__142;
  assign wide_x__59 = {2'h1, x_fraction__235, 3'h0};
  assign result_sign__240 = x_sign__92 & prod_sign__46 & concat_165662[0] | ~prod_sign__46 & concat_165662[1] | prod_sign__46 & concat_165662[2];
  assign x_fraction__380 = sum__50[8] ? result_fraction__294 : result_fraction__300;
  assign dropped__50 = sub_165668 >= 8'h1c ? 28'h000_0000 : wide_y__100 << sub_165668;
  assign result_sign__241 = is_operand_inf__47 ? ~has_pos_inf__47 : result_sign__239;
  assign wide_x__97 = {2'h1, x_fraction__379, 3'h0};
  assign result_sign__337 = x_sign__128 & prod_sign__64 & concat_165676[0] | ~prod_sign__64 & concat_165676[1] | prod_sign__64 & concat_165676[2];
  assign x_fraction__524 = sum__69[8] ? result_fraction__411 : result_fraction__417;
  assign dropped__69 = sub_165682 >= 8'h1c ? 28'h000_0000 : wide_y__138 << sub_165682;
  assign x_sign__129 = array_index_164412[31:31];
  assign result_sign__338 = is_operand_inf__66 ? ~has_pos_inf__66 : result_sign__336;
  assign wide_x__135 = {2'h1, x_fraction__523, 3'h0};
  assign result_sign__24 = is_operand_inf__5 ? ~has_pos_inf__5 : result_sign__23;
  assign wide_x__11 = {2'h1, x_fraction__46, 3'h0};
  assign result_sign__69 = ~is_result_nan__27 & result_sign__68;
  assign wide_x__29 = wide_x__28 & {28{x_bexp__118 != x_bexp__752}};
  assign result_sign__145 = is_operand_inf__29 ? ~has_pos_inf__29 : result_sign__143;
  assign wide_x__60 = {2'h1, x_fraction__236, 3'h0};
  assign result_sign__150 = x_bexp__461 != high_exp__482 & x_sign__117;
  assign result_sign__146 = ~is_result_nan__58 & result_sign__144;
  assign wide_x__61 = wide_x__59 & {28{x_bexp__235 != x_bexp__753}};
  assign result_sign__242 = is_operand_inf__48 ? ~has_pos_inf__48 : result_sign__240;
  assign wide_x__98 = {2'h1, x_fraction__380, 3'h0};
  assign result_sign__243 = ~is_result_nan__97 & result_sign__241;
  assign wide_x__99 = wide_x__97 & {28{x_bexp__379 != x_bexp__754}};
  assign result_sign__339 = is_operand_inf__67 ? ~has_pos_inf__67 : result_sign__337;
  assign wide_x__136 = {2'h1, x_fraction__524, 3'h0};
  assign result_sign__344 = x_bexp__510 != high_exp__489 & x_sign__129;
  assign result_sign__340 = ~is_result_nan__136 & result_sign__338;
  assign wide_x__137 = wide_x__135 & {28{x_bexp__523 != x_bexp__755}};
  assign result_sign__25 = ~is_result_nan__10 & result_sign__24;
  assign wide_x__12 = wide_x__11 & {28{x_bexp__46 != x_bexp__756}};
  assign x_sign__30 = sum__14[8] ? result_sign__69 : result_sign__305;
  assign prod_sign__14 = sum__14[8] ? result_sign__305 : result_sign__69;
  assign neg_165796 = -wide_x__29;
  assign sticky__44 = {27'h000_0000, dropped__14[27:3] != 25'h000_0000};
  assign result_sign__147 = ~is_result_nan__59 & result_sign__145;
  assign wide_x__62 = wide_x__60 & {28{x_bexp__236 != x_bexp__757}};
  assign x_sign__59 = sum__30[8] ? result_sign__146 : result_sign__150;
  assign prod_sign__29 = sum__30[8] ? result_sign__150 : result_sign__146;
  assign neg_165805 = -wide_x__61;
  assign sticky__94 = {27'h000_0000, dropped__30[27:3] != 25'h000_0000};
  assign result_sign__248 = ~(is_result_nan__134 & ne_165126) & x_sign__125;
  assign result_sign__244 = ~is_result_nan__98 & result_sign__242;
  assign wide_x__100 = wide_x__98 & {28{x_bexp__380 != x_bexp__758}};
  assign x_sign__95 = sum__49[8] ? result_sign__243 : result_sign__334;
  assign prod_sign__47 = sum__49[8] ? result_sign__334 : result_sign__243;
  assign neg_165815 = -wide_x__99;
  assign sticky__153 = {27'h000_0000, dropped__49[27:3] != 25'h000_0000};
  assign result_sign__345 = ~(is_result_nan__138 & ne_165140) & x_sign__129;
  assign result_sign__341 = ~is_result_nan__137 & result_sign__339;
  assign wide_x__138 = wide_x__136 & {28{x_bexp__524 != x_bexp__759}};
  assign x_sign__131 = sum__68[8] ? result_sign__340 : result_sign__344;
  assign prod_sign__65 = sum__68[8] ? result_sign__344 : result_sign__340;
  assign neg_165825 = -wide_x__137;
  assign sticky__212 = {27'h000_0000, dropped__68[27:3] != 25'h000_0000};
  assign x_sign__12 = sum__6[8] ? result_sign__25 : result_sign__218;
  assign prod_sign__6 = sum__6[8] ? result_sign__218 : result_sign__25;
  assign neg_165830 = -wide_x__12;
  assign sticky__18 = {27'h000_0000, dropped__6[27:3] != 25'h000_0000};
  assign xddend_y__14 = (x_bexpbs_difference__15 >= 8'h1c ? 28'h000_0000 : wide_y__29 >> x_bexpbs_difference__15) | sticky__44;
  assign x_sign__60 = sum__31[8] ? result_sign__147 : result_sign__315;
  assign prod_sign__30 = sum__31[8] ? result_sign__315 : result_sign__147;
  assign neg_165839 = -wide_x__62;
  assign sticky__95 = {27'h000_0000, dropped__31[27:3] != 25'h000_0000};
  assign xddend_y__29 = (x_bexpbs_difference__29 >= 8'h1c ? 28'h000_0000 : wide_y__61 >> x_bexpbs_difference__29) | sticky__94;
  assign x_sign__96 = sum__50[8] ? result_sign__244 : result_sign__248;
  assign prod_sign__48 = sum__50[8] ? result_sign__248 : result_sign__244;
  assign neg_165848 = -wide_x__100;
  assign sticky__154 = {27'h000_0000, dropped__50[27:3] != 25'h000_0000};
  assign xddend_y__47 = (x_bexpbs_difference__47 >= 8'h1c ? 28'h000_0000 : wide_y__99 >> x_bexpbs_difference__47) | sticky__153;
  assign x_sign__132 = sum__69[8] ? result_sign__341 : result_sign__345;
  assign prod_sign__66 = sum__69[8] ? result_sign__345 : result_sign__341;
  assign neg_165857 = -wide_x__138;
  assign sticky__213 = {27'h000_0000, dropped__69[27:3] != 25'h000_0000};
  assign xddend_y__65 = (x_bexpbs_difference__65 >= 8'h1c ? 28'h000_0000 : wide_y__137 >> x_bexpbs_difference__65) | sticky__212;
  assign xddend_y__6 = (x_bexpbs_difference__6 >= 8'h1c ? 28'h000_0000 : wide_y__12 >> x_bexpbs_difference__6) | sticky__18;
  assign sel_165868 = x_sign__30 ^ prod_sign__14 ? neg_165796[27:3] : wide_x__29[27:3];
  assign result_sign__1034 = 1'h0;
  assign xddend_y__30 = (x_bexpbs_difference__30 >= 8'h1c ? 28'h000_0000 : wide_y__62 >> x_bexpbs_difference__30) | sticky__95;
  assign sel_165875 = x_sign__59 ^ prod_sign__29 ? neg_165805[27:3] : wide_x__61[27:3];
  assign result_sign__1035 = 1'h0;
  assign xddend_y__48 = (x_bexpbs_difference__48 >= 8'h1c ? 28'h000_0000 : wide_y__100 >> x_bexpbs_difference__48) | sticky__154;
  assign sel_165882 = x_sign__95 ^ prod_sign__47 ? neg_165815[27:3] : wide_x__99[27:3];
  assign result_sign__1036 = 1'h0;
  assign xddend_y__66 = (x_bexpbs_difference__66 >= 8'h1c ? 28'h000_0000 : wide_y__138 >> x_bexpbs_difference__66) | sticky__213;
  assign sel_165889 = x_sign__131 ^ prod_sign__65 ? neg_165825[27:3] : wide_x__137[27:3];
  assign result_sign__1037 = 1'h0;
  assign sel_165892 = x_sign__12 ^ prod_sign__6 ? neg_165830[27:3] : wide_x__12[27:3];
  assign result_sign__1038 = 1'h0;
  assign sel_165897 = x_sign__60 ^ prod_sign__30 ? neg_165839[27:3] : wide_x__62[27:3];
  assign result_sign__1039 = 1'h0;
  assign sel_165902 = x_sign__96 ^ prod_sign__48 ? neg_165848[27:3] : wide_x__100[27:3];
  assign result_sign__1040 = 1'h0;
  assign sel_165907 = x_sign__132 ^ prod_sign__66 ? neg_165857[27:3] : wide_x__138[27:3];
  assign result_sign__1041 = 1'h0;
  assign add_165914 = {{1{sel_165868[24]}}, sel_165868} + {result_sign__1034, xddend_y__14[27:3]};
  assign add_165917 = {{1{sel_165875[24]}}, sel_165875} + {result_sign__1035, xddend_y__29[27:3]};
  assign add_165920 = {{1{sel_165882[24]}}, sel_165882} + {result_sign__1036, xddend_y__47[27:3]};
  assign add_165923 = {{1{sel_165889[24]}}, sel_165889} + {result_sign__1037, xddend_y__65[27:3]};
  assign add_165924 = {{1{sel_165892[24]}}, sel_165892} + {result_sign__1038, xddend_y__6[27:3]};
  assign add_165927 = {{1{sel_165897[24]}}, sel_165897} + {result_sign__1039, xddend_y__30[27:3]};
  assign add_165930 = {{1{sel_165902[24]}}, sel_165902} + {result_sign__1040, xddend_y__48[27:3]};
  assign add_165933 = {{1{sel_165907[24]}}, sel_165907} + {result_sign__1041, xddend_y__66[27:3]};
  assign concat_165938 = {add_165914[24:0], xddend_y__14[2:0]};
  assign concat_165941 = {add_165917[24:0], xddend_y__29[2:0]};
  assign concat_165944 = {add_165920[24:0], xddend_y__47[2:0]};
  assign concat_165947 = {add_165923[24:0], xddend_y__65[2:0]};
  assign concat_165948 = {add_165924[24:0], xddend_y__6[2:0]};
  assign concat_165951 = {add_165927[24:0], xddend_y__30[2:0]};
  assign concat_165954 = {add_165930[24:0], xddend_y__48[2:0]};
  assign concat_165957 = {add_165933[24:0], xddend_y__66[2:0]};
  assign xbs_fraction__14 = add_165914[25] ? -concat_165938 : concat_165938;
  assign xbs_fraction__29 = add_165917[25] ? -concat_165941 : concat_165941;
  assign xbs_fraction__47 = add_165920[25] ? -concat_165944 : concat_165944;
  assign xbs_fraction__65 = add_165923[25] ? -concat_165947 : concat_165947;
  assign xbs_fraction__6 = add_165924[25] ? -concat_165948 : concat_165948;
  assign reverse_165973 = {xbs_fraction__14[0], xbs_fraction__14[1], xbs_fraction__14[2], xbs_fraction__14[3], xbs_fraction__14[4], xbs_fraction__14[5], xbs_fraction__14[6], xbs_fraction__14[7], xbs_fraction__14[8], xbs_fraction__14[9], xbs_fraction__14[10], xbs_fraction__14[11], xbs_fraction__14[12], xbs_fraction__14[13], xbs_fraction__14[14], xbs_fraction__14[15], xbs_fraction__14[16], xbs_fraction__14[17], xbs_fraction__14[18], xbs_fraction__14[19], xbs_fraction__14[20], xbs_fraction__14[21], xbs_fraction__14[22], xbs_fraction__14[23], xbs_fraction__14[24], xbs_fraction__14[25], xbs_fraction__14[26], xbs_fraction__14[27]};
  assign xbs_fraction__30 = add_165927[25] ? -concat_165951 : concat_165951;
  assign reverse_165975 = {xbs_fraction__29[0], xbs_fraction__29[1], xbs_fraction__29[2], xbs_fraction__29[3], xbs_fraction__29[4], xbs_fraction__29[5], xbs_fraction__29[6], xbs_fraction__29[7], xbs_fraction__29[8], xbs_fraction__29[9], xbs_fraction__29[10], xbs_fraction__29[11], xbs_fraction__29[12], xbs_fraction__29[13], xbs_fraction__29[14], xbs_fraction__29[15], xbs_fraction__29[16], xbs_fraction__29[17], xbs_fraction__29[18], xbs_fraction__29[19], xbs_fraction__29[20], xbs_fraction__29[21], xbs_fraction__29[22], xbs_fraction__29[23], xbs_fraction__29[24], xbs_fraction__29[25], xbs_fraction__29[26], xbs_fraction__29[27]};
  assign xbs_fraction__48 = add_165930[25] ? -concat_165954 : concat_165954;
  assign reverse_165977 = {xbs_fraction__47[0], xbs_fraction__47[1], xbs_fraction__47[2], xbs_fraction__47[3], xbs_fraction__47[4], xbs_fraction__47[5], xbs_fraction__47[6], xbs_fraction__47[7], xbs_fraction__47[8], xbs_fraction__47[9], xbs_fraction__47[10], xbs_fraction__47[11], xbs_fraction__47[12], xbs_fraction__47[13], xbs_fraction__47[14], xbs_fraction__47[15], xbs_fraction__47[16], xbs_fraction__47[17], xbs_fraction__47[18], xbs_fraction__47[19], xbs_fraction__47[20], xbs_fraction__47[21], xbs_fraction__47[22], xbs_fraction__47[23], xbs_fraction__47[24], xbs_fraction__47[25], xbs_fraction__47[26], xbs_fraction__47[27]};
  assign xbs_fraction__66 = add_165933[25] ? -concat_165957 : concat_165957;
  assign reverse_165979 = {xbs_fraction__65[0], xbs_fraction__65[1], xbs_fraction__65[2], xbs_fraction__65[3], xbs_fraction__65[4], xbs_fraction__65[5], xbs_fraction__65[6], xbs_fraction__65[7], xbs_fraction__65[8], xbs_fraction__65[9], xbs_fraction__65[10], xbs_fraction__65[11], xbs_fraction__65[12], xbs_fraction__65[13], xbs_fraction__65[14], xbs_fraction__65[15], xbs_fraction__65[16], xbs_fraction__65[17], xbs_fraction__65[18], xbs_fraction__65[19], xbs_fraction__65[20], xbs_fraction__65[21], xbs_fraction__65[22], xbs_fraction__65[23], xbs_fraction__65[24], xbs_fraction__65[25], xbs_fraction__65[26], xbs_fraction__65[27]};
  assign reverse_165980 = {xbs_fraction__6[0], xbs_fraction__6[1], xbs_fraction__6[2], xbs_fraction__6[3], xbs_fraction__6[4], xbs_fraction__6[5], xbs_fraction__6[6], xbs_fraction__6[7], xbs_fraction__6[8], xbs_fraction__6[9], xbs_fraction__6[10], xbs_fraction__6[11], xbs_fraction__6[12], xbs_fraction__6[13], xbs_fraction__6[14], xbs_fraction__6[15], xbs_fraction__6[16], xbs_fraction__6[17], xbs_fraction__6[18], xbs_fraction__6[19], xbs_fraction__6[20], xbs_fraction__6[21], xbs_fraction__6[22], xbs_fraction__6[23], xbs_fraction__6[24], xbs_fraction__6[25], xbs_fraction__6[26], xbs_fraction__6[27]};
  assign one_hot_165981 = {reverse_165973[27:0] == 28'h000_0000, reverse_165973[27] && reverse_165973[26:0] == 27'h000_0000, reverse_165973[26] && reverse_165973[25:0] == 26'h000_0000, reverse_165973[25] && reverse_165973[24:0] == 25'h000_0000, reverse_165973[24] && reverse_165973[23:0] == 24'h00_0000, reverse_165973[23] && reverse_165973[22:0] == 23'h00_0000, reverse_165973[22] && reverse_165973[21:0] == 22'h00_0000, reverse_165973[21] && reverse_165973[20:0] == 21'h00_0000, reverse_165973[20] && reverse_165973[19:0] == 20'h0_0000, reverse_165973[19] && reverse_165973[18:0] == 19'h0_0000, reverse_165973[18] && reverse_165973[17:0] == 18'h0_0000, reverse_165973[17] && reverse_165973[16:0] == 17'h0_0000, reverse_165973[16] && reverse_165973[15:0] == 16'h0000, reverse_165973[15] && reverse_165973[14:0] == 15'h0000, reverse_165973[14] && reverse_165973[13:0] == 14'h0000, reverse_165973[13] && reverse_165973[12:0] == 13'h0000, reverse_165973[12] && reverse_165973[11:0] == 12'h000, reverse_165973[11] && reverse_165973[10:0] == 11'h000, reverse_165973[10] && reverse_165973[9:0] == 10'h000, reverse_165973[9] && reverse_165973[8:0] == 9'h000, reverse_165973[8] && reverse_165973[7:0] == 8'h00, reverse_165973[7] && reverse_165973[6:0] == 7'h00, reverse_165973[6] && reverse_165973[5:0] == 6'h00, reverse_165973[5] && reverse_165973[4:0] == 5'h00, reverse_165973[4] && reverse_165973[3:0] == 4'h0, reverse_165973[3] && reverse_165973[2:0] == 3'h0, reverse_165973[2] && reverse_165973[1:0] == 2'h0, reverse_165973[1] && !reverse_165973[0], reverse_165973[0]};
  assign reverse_165982 = {xbs_fraction__30[0], xbs_fraction__30[1], xbs_fraction__30[2], xbs_fraction__30[3], xbs_fraction__30[4], xbs_fraction__30[5], xbs_fraction__30[6], xbs_fraction__30[7], xbs_fraction__30[8], xbs_fraction__30[9], xbs_fraction__30[10], xbs_fraction__30[11], xbs_fraction__30[12], xbs_fraction__30[13], xbs_fraction__30[14], xbs_fraction__30[15], xbs_fraction__30[16], xbs_fraction__30[17], xbs_fraction__30[18], xbs_fraction__30[19], xbs_fraction__30[20], xbs_fraction__30[21], xbs_fraction__30[22], xbs_fraction__30[23], xbs_fraction__30[24], xbs_fraction__30[25], xbs_fraction__30[26], xbs_fraction__30[27]};
  assign one_hot_165983 = {reverse_165975[27:0] == 28'h000_0000, reverse_165975[27] && reverse_165975[26:0] == 27'h000_0000, reverse_165975[26] && reverse_165975[25:0] == 26'h000_0000, reverse_165975[25] && reverse_165975[24:0] == 25'h000_0000, reverse_165975[24] && reverse_165975[23:0] == 24'h00_0000, reverse_165975[23] && reverse_165975[22:0] == 23'h00_0000, reverse_165975[22] && reverse_165975[21:0] == 22'h00_0000, reverse_165975[21] && reverse_165975[20:0] == 21'h00_0000, reverse_165975[20] && reverse_165975[19:0] == 20'h0_0000, reverse_165975[19] && reverse_165975[18:0] == 19'h0_0000, reverse_165975[18] && reverse_165975[17:0] == 18'h0_0000, reverse_165975[17] && reverse_165975[16:0] == 17'h0_0000, reverse_165975[16] && reverse_165975[15:0] == 16'h0000, reverse_165975[15] && reverse_165975[14:0] == 15'h0000, reverse_165975[14] && reverse_165975[13:0] == 14'h0000, reverse_165975[13] && reverse_165975[12:0] == 13'h0000, reverse_165975[12] && reverse_165975[11:0] == 12'h000, reverse_165975[11] && reverse_165975[10:0] == 11'h000, reverse_165975[10] && reverse_165975[9:0] == 10'h000, reverse_165975[9] && reverse_165975[8:0] == 9'h000, reverse_165975[8] && reverse_165975[7:0] == 8'h00, reverse_165975[7] && reverse_165975[6:0] == 7'h00, reverse_165975[6] && reverse_165975[5:0] == 6'h00, reverse_165975[5] && reverse_165975[4:0] == 5'h00, reverse_165975[4] && reverse_165975[3:0] == 4'h0, reverse_165975[3] && reverse_165975[2:0] == 3'h0, reverse_165975[2] && reverse_165975[1:0] == 2'h0, reverse_165975[1] && !reverse_165975[0], reverse_165975[0]};
  assign reverse_165984 = {xbs_fraction__48[0], xbs_fraction__48[1], xbs_fraction__48[2], xbs_fraction__48[3], xbs_fraction__48[4], xbs_fraction__48[5], xbs_fraction__48[6], xbs_fraction__48[7], xbs_fraction__48[8], xbs_fraction__48[9], xbs_fraction__48[10], xbs_fraction__48[11], xbs_fraction__48[12], xbs_fraction__48[13], xbs_fraction__48[14], xbs_fraction__48[15], xbs_fraction__48[16], xbs_fraction__48[17], xbs_fraction__48[18], xbs_fraction__48[19], xbs_fraction__48[20], xbs_fraction__48[21], xbs_fraction__48[22], xbs_fraction__48[23], xbs_fraction__48[24], xbs_fraction__48[25], xbs_fraction__48[26], xbs_fraction__48[27]};
  assign one_hot_165985 = {reverse_165977[27:0] == 28'h000_0000, reverse_165977[27] && reverse_165977[26:0] == 27'h000_0000, reverse_165977[26] && reverse_165977[25:0] == 26'h000_0000, reverse_165977[25] && reverse_165977[24:0] == 25'h000_0000, reverse_165977[24] && reverse_165977[23:0] == 24'h00_0000, reverse_165977[23] && reverse_165977[22:0] == 23'h00_0000, reverse_165977[22] && reverse_165977[21:0] == 22'h00_0000, reverse_165977[21] && reverse_165977[20:0] == 21'h00_0000, reverse_165977[20] && reverse_165977[19:0] == 20'h0_0000, reverse_165977[19] && reverse_165977[18:0] == 19'h0_0000, reverse_165977[18] && reverse_165977[17:0] == 18'h0_0000, reverse_165977[17] && reverse_165977[16:0] == 17'h0_0000, reverse_165977[16] && reverse_165977[15:0] == 16'h0000, reverse_165977[15] && reverse_165977[14:0] == 15'h0000, reverse_165977[14] && reverse_165977[13:0] == 14'h0000, reverse_165977[13] && reverse_165977[12:0] == 13'h0000, reverse_165977[12] && reverse_165977[11:0] == 12'h000, reverse_165977[11] && reverse_165977[10:0] == 11'h000, reverse_165977[10] && reverse_165977[9:0] == 10'h000, reverse_165977[9] && reverse_165977[8:0] == 9'h000, reverse_165977[8] && reverse_165977[7:0] == 8'h00, reverse_165977[7] && reverse_165977[6:0] == 7'h00, reverse_165977[6] && reverse_165977[5:0] == 6'h00, reverse_165977[5] && reverse_165977[4:0] == 5'h00, reverse_165977[4] && reverse_165977[3:0] == 4'h0, reverse_165977[3] && reverse_165977[2:0] == 3'h0, reverse_165977[2] && reverse_165977[1:0] == 2'h0, reverse_165977[1] && !reverse_165977[0], reverse_165977[0]};
  assign reverse_165986 = {xbs_fraction__66[0], xbs_fraction__66[1], xbs_fraction__66[2], xbs_fraction__66[3], xbs_fraction__66[4], xbs_fraction__66[5], xbs_fraction__66[6], xbs_fraction__66[7], xbs_fraction__66[8], xbs_fraction__66[9], xbs_fraction__66[10], xbs_fraction__66[11], xbs_fraction__66[12], xbs_fraction__66[13], xbs_fraction__66[14], xbs_fraction__66[15], xbs_fraction__66[16], xbs_fraction__66[17], xbs_fraction__66[18], xbs_fraction__66[19], xbs_fraction__66[20], xbs_fraction__66[21], xbs_fraction__66[22], xbs_fraction__66[23], xbs_fraction__66[24], xbs_fraction__66[25], xbs_fraction__66[26], xbs_fraction__66[27]};
  assign one_hot_165987 = {reverse_165979[27:0] == 28'h000_0000, reverse_165979[27] && reverse_165979[26:0] == 27'h000_0000, reverse_165979[26] && reverse_165979[25:0] == 26'h000_0000, reverse_165979[25] && reverse_165979[24:0] == 25'h000_0000, reverse_165979[24] && reverse_165979[23:0] == 24'h00_0000, reverse_165979[23] && reverse_165979[22:0] == 23'h00_0000, reverse_165979[22] && reverse_165979[21:0] == 22'h00_0000, reverse_165979[21] && reverse_165979[20:0] == 21'h00_0000, reverse_165979[20] && reverse_165979[19:0] == 20'h0_0000, reverse_165979[19] && reverse_165979[18:0] == 19'h0_0000, reverse_165979[18] && reverse_165979[17:0] == 18'h0_0000, reverse_165979[17] && reverse_165979[16:0] == 17'h0_0000, reverse_165979[16] && reverse_165979[15:0] == 16'h0000, reverse_165979[15] && reverse_165979[14:0] == 15'h0000, reverse_165979[14] && reverse_165979[13:0] == 14'h0000, reverse_165979[13] && reverse_165979[12:0] == 13'h0000, reverse_165979[12] && reverse_165979[11:0] == 12'h000, reverse_165979[11] && reverse_165979[10:0] == 11'h000, reverse_165979[10] && reverse_165979[9:0] == 10'h000, reverse_165979[9] && reverse_165979[8:0] == 9'h000, reverse_165979[8] && reverse_165979[7:0] == 8'h00, reverse_165979[7] && reverse_165979[6:0] == 7'h00, reverse_165979[6] && reverse_165979[5:0] == 6'h00, reverse_165979[5] && reverse_165979[4:0] == 5'h00, reverse_165979[4] && reverse_165979[3:0] == 4'h0, reverse_165979[3] && reverse_165979[2:0] == 3'h0, reverse_165979[2] && reverse_165979[1:0] == 2'h0, reverse_165979[1] && !reverse_165979[0], reverse_165979[0]};
  assign one_hot_165988 = {reverse_165980[27:0] == 28'h000_0000, reverse_165980[27] && reverse_165980[26:0] == 27'h000_0000, reverse_165980[26] && reverse_165980[25:0] == 26'h000_0000, reverse_165980[25] && reverse_165980[24:0] == 25'h000_0000, reverse_165980[24] && reverse_165980[23:0] == 24'h00_0000, reverse_165980[23] && reverse_165980[22:0] == 23'h00_0000, reverse_165980[22] && reverse_165980[21:0] == 22'h00_0000, reverse_165980[21] && reverse_165980[20:0] == 21'h00_0000, reverse_165980[20] && reverse_165980[19:0] == 20'h0_0000, reverse_165980[19] && reverse_165980[18:0] == 19'h0_0000, reverse_165980[18] && reverse_165980[17:0] == 18'h0_0000, reverse_165980[17] && reverse_165980[16:0] == 17'h0_0000, reverse_165980[16] && reverse_165980[15:0] == 16'h0000, reverse_165980[15] && reverse_165980[14:0] == 15'h0000, reverse_165980[14] && reverse_165980[13:0] == 14'h0000, reverse_165980[13] && reverse_165980[12:0] == 13'h0000, reverse_165980[12] && reverse_165980[11:0] == 12'h000, reverse_165980[11] && reverse_165980[10:0] == 11'h000, reverse_165980[10] && reverse_165980[9:0] == 10'h000, reverse_165980[9] && reverse_165980[8:0] == 9'h000, reverse_165980[8] && reverse_165980[7:0] == 8'h00, reverse_165980[7] && reverse_165980[6:0] == 7'h00, reverse_165980[6] && reverse_165980[5:0] == 6'h00, reverse_165980[5] && reverse_165980[4:0] == 5'h00, reverse_165980[4] && reverse_165980[3:0] == 4'h0, reverse_165980[3] && reverse_165980[2:0] == 3'h0, reverse_165980[2] && reverse_165980[1:0] == 2'h0, reverse_165980[1] && !reverse_165980[0], reverse_165980[0]};
  assign encode_165989 = {one_hot_165981[16] | one_hot_165981[17] | one_hot_165981[18] | one_hot_165981[19] | one_hot_165981[20] | one_hot_165981[21] | one_hot_165981[22] | one_hot_165981[23] | one_hot_165981[24] | one_hot_165981[25] | one_hot_165981[26] | one_hot_165981[27] | one_hot_165981[28], one_hot_165981[8] | one_hot_165981[9] | one_hot_165981[10] | one_hot_165981[11] | one_hot_165981[12] | one_hot_165981[13] | one_hot_165981[14] | one_hot_165981[15] | one_hot_165981[24] | one_hot_165981[25] | one_hot_165981[26] | one_hot_165981[27] | one_hot_165981[28], one_hot_165981[4] | one_hot_165981[5] | one_hot_165981[6] | one_hot_165981[7] | one_hot_165981[12] | one_hot_165981[13] | one_hot_165981[14] | one_hot_165981[15] | one_hot_165981[20] | one_hot_165981[21] | one_hot_165981[22] | one_hot_165981[23] | one_hot_165981[28], one_hot_165981[2] | one_hot_165981[3] | one_hot_165981[6] | one_hot_165981[7] | one_hot_165981[10] | one_hot_165981[11] | one_hot_165981[14] | one_hot_165981[15] | one_hot_165981[18] | one_hot_165981[19] | one_hot_165981[22] | one_hot_165981[23] | one_hot_165981[26] | one_hot_165981[27], one_hot_165981[1] | one_hot_165981[3] | one_hot_165981[5] | one_hot_165981[7] | one_hot_165981[9] | one_hot_165981[11] | one_hot_165981[13] | one_hot_165981[15] | one_hot_165981[17] | one_hot_165981[19] | one_hot_165981[21] | one_hot_165981[23] | one_hot_165981[25] | one_hot_165981[27]};
  assign one_hot_165990 = {reverse_165982[27:0] == 28'h000_0000, reverse_165982[27] && reverse_165982[26:0] == 27'h000_0000, reverse_165982[26] && reverse_165982[25:0] == 26'h000_0000, reverse_165982[25] && reverse_165982[24:0] == 25'h000_0000, reverse_165982[24] && reverse_165982[23:0] == 24'h00_0000, reverse_165982[23] && reverse_165982[22:0] == 23'h00_0000, reverse_165982[22] && reverse_165982[21:0] == 22'h00_0000, reverse_165982[21] && reverse_165982[20:0] == 21'h00_0000, reverse_165982[20] && reverse_165982[19:0] == 20'h0_0000, reverse_165982[19] && reverse_165982[18:0] == 19'h0_0000, reverse_165982[18] && reverse_165982[17:0] == 18'h0_0000, reverse_165982[17] && reverse_165982[16:0] == 17'h0_0000, reverse_165982[16] && reverse_165982[15:0] == 16'h0000, reverse_165982[15] && reverse_165982[14:0] == 15'h0000, reverse_165982[14] && reverse_165982[13:0] == 14'h0000, reverse_165982[13] && reverse_165982[12:0] == 13'h0000, reverse_165982[12] && reverse_165982[11:0] == 12'h000, reverse_165982[11] && reverse_165982[10:0] == 11'h000, reverse_165982[10] && reverse_165982[9:0] == 10'h000, reverse_165982[9] && reverse_165982[8:0] == 9'h000, reverse_165982[8] && reverse_165982[7:0] == 8'h00, reverse_165982[7] && reverse_165982[6:0] == 7'h00, reverse_165982[6] && reverse_165982[5:0] == 6'h00, reverse_165982[5] && reverse_165982[4:0] == 5'h00, reverse_165982[4] && reverse_165982[3:0] == 4'h0, reverse_165982[3] && reverse_165982[2:0] == 3'h0, reverse_165982[2] && reverse_165982[1:0] == 2'h0, reverse_165982[1] && !reverse_165982[0], reverse_165982[0]};
  assign encode_165991 = {one_hot_165983[16] | one_hot_165983[17] | one_hot_165983[18] | one_hot_165983[19] | one_hot_165983[20] | one_hot_165983[21] | one_hot_165983[22] | one_hot_165983[23] | one_hot_165983[24] | one_hot_165983[25] | one_hot_165983[26] | one_hot_165983[27] | one_hot_165983[28], one_hot_165983[8] | one_hot_165983[9] | one_hot_165983[10] | one_hot_165983[11] | one_hot_165983[12] | one_hot_165983[13] | one_hot_165983[14] | one_hot_165983[15] | one_hot_165983[24] | one_hot_165983[25] | one_hot_165983[26] | one_hot_165983[27] | one_hot_165983[28], one_hot_165983[4] | one_hot_165983[5] | one_hot_165983[6] | one_hot_165983[7] | one_hot_165983[12] | one_hot_165983[13] | one_hot_165983[14] | one_hot_165983[15] | one_hot_165983[20] | one_hot_165983[21] | one_hot_165983[22] | one_hot_165983[23] | one_hot_165983[28], one_hot_165983[2] | one_hot_165983[3] | one_hot_165983[6] | one_hot_165983[7] | one_hot_165983[10] | one_hot_165983[11] | one_hot_165983[14] | one_hot_165983[15] | one_hot_165983[18] | one_hot_165983[19] | one_hot_165983[22] | one_hot_165983[23] | one_hot_165983[26] | one_hot_165983[27], one_hot_165983[1] | one_hot_165983[3] | one_hot_165983[5] | one_hot_165983[7] | one_hot_165983[9] | one_hot_165983[11] | one_hot_165983[13] | one_hot_165983[15] | one_hot_165983[17] | one_hot_165983[19] | one_hot_165983[21] | one_hot_165983[23] | one_hot_165983[25] | one_hot_165983[27]};
  assign one_hot_165992 = {reverse_165984[27:0] == 28'h000_0000, reverse_165984[27] && reverse_165984[26:0] == 27'h000_0000, reverse_165984[26] && reverse_165984[25:0] == 26'h000_0000, reverse_165984[25] && reverse_165984[24:0] == 25'h000_0000, reverse_165984[24] && reverse_165984[23:0] == 24'h00_0000, reverse_165984[23] && reverse_165984[22:0] == 23'h00_0000, reverse_165984[22] && reverse_165984[21:0] == 22'h00_0000, reverse_165984[21] && reverse_165984[20:0] == 21'h00_0000, reverse_165984[20] && reverse_165984[19:0] == 20'h0_0000, reverse_165984[19] && reverse_165984[18:0] == 19'h0_0000, reverse_165984[18] && reverse_165984[17:0] == 18'h0_0000, reverse_165984[17] && reverse_165984[16:0] == 17'h0_0000, reverse_165984[16] && reverse_165984[15:0] == 16'h0000, reverse_165984[15] && reverse_165984[14:0] == 15'h0000, reverse_165984[14] && reverse_165984[13:0] == 14'h0000, reverse_165984[13] && reverse_165984[12:0] == 13'h0000, reverse_165984[12] && reverse_165984[11:0] == 12'h000, reverse_165984[11] && reverse_165984[10:0] == 11'h000, reverse_165984[10] && reverse_165984[9:0] == 10'h000, reverse_165984[9] && reverse_165984[8:0] == 9'h000, reverse_165984[8] && reverse_165984[7:0] == 8'h00, reverse_165984[7] && reverse_165984[6:0] == 7'h00, reverse_165984[6] && reverse_165984[5:0] == 6'h00, reverse_165984[5] && reverse_165984[4:0] == 5'h00, reverse_165984[4] && reverse_165984[3:0] == 4'h0, reverse_165984[3] && reverse_165984[2:0] == 3'h0, reverse_165984[2] && reverse_165984[1:0] == 2'h0, reverse_165984[1] && !reverse_165984[0], reverse_165984[0]};
  assign encode_165993 = {one_hot_165985[16] | one_hot_165985[17] | one_hot_165985[18] | one_hot_165985[19] | one_hot_165985[20] | one_hot_165985[21] | one_hot_165985[22] | one_hot_165985[23] | one_hot_165985[24] | one_hot_165985[25] | one_hot_165985[26] | one_hot_165985[27] | one_hot_165985[28], one_hot_165985[8] | one_hot_165985[9] | one_hot_165985[10] | one_hot_165985[11] | one_hot_165985[12] | one_hot_165985[13] | one_hot_165985[14] | one_hot_165985[15] | one_hot_165985[24] | one_hot_165985[25] | one_hot_165985[26] | one_hot_165985[27] | one_hot_165985[28], one_hot_165985[4] | one_hot_165985[5] | one_hot_165985[6] | one_hot_165985[7] | one_hot_165985[12] | one_hot_165985[13] | one_hot_165985[14] | one_hot_165985[15] | one_hot_165985[20] | one_hot_165985[21] | one_hot_165985[22] | one_hot_165985[23] | one_hot_165985[28], one_hot_165985[2] | one_hot_165985[3] | one_hot_165985[6] | one_hot_165985[7] | one_hot_165985[10] | one_hot_165985[11] | one_hot_165985[14] | one_hot_165985[15] | one_hot_165985[18] | one_hot_165985[19] | one_hot_165985[22] | one_hot_165985[23] | one_hot_165985[26] | one_hot_165985[27], one_hot_165985[1] | one_hot_165985[3] | one_hot_165985[5] | one_hot_165985[7] | one_hot_165985[9] | one_hot_165985[11] | one_hot_165985[13] | one_hot_165985[15] | one_hot_165985[17] | one_hot_165985[19] | one_hot_165985[21] | one_hot_165985[23] | one_hot_165985[25] | one_hot_165985[27]};
  assign one_hot_165994 = {reverse_165986[27:0] == 28'h000_0000, reverse_165986[27] && reverse_165986[26:0] == 27'h000_0000, reverse_165986[26] && reverse_165986[25:0] == 26'h000_0000, reverse_165986[25] && reverse_165986[24:0] == 25'h000_0000, reverse_165986[24] && reverse_165986[23:0] == 24'h00_0000, reverse_165986[23] && reverse_165986[22:0] == 23'h00_0000, reverse_165986[22] && reverse_165986[21:0] == 22'h00_0000, reverse_165986[21] && reverse_165986[20:0] == 21'h00_0000, reverse_165986[20] && reverse_165986[19:0] == 20'h0_0000, reverse_165986[19] && reverse_165986[18:0] == 19'h0_0000, reverse_165986[18] && reverse_165986[17:0] == 18'h0_0000, reverse_165986[17] && reverse_165986[16:0] == 17'h0_0000, reverse_165986[16] && reverse_165986[15:0] == 16'h0000, reverse_165986[15] && reverse_165986[14:0] == 15'h0000, reverse_165986[14] && reverse_165986[13:0] == 14'h0000, reverse_165986[13] && reverse_165986[12:0] == 13'h0000, reverse_165986[12] && reverse_165986[11:0] == 12'h000, reverse_165986[11] && reverse_165986[10:0] == 11'h000, reverse_165986[10] && reverse_165986[9:0] == 10'h000, reverse_165986[9] && reverse_165986[8:0] == 9'h000, reverse_165986[8] && reverse_165986[7:0] == 8'h00, reverse_165986[7] && reverse_165986[6:0] == 7'h00, reverse_165986[6] && reverse_165986[5:0] == 6'h00, reverse_165986[5] && reverse_165986[4:0] == 5'h00, reverse_165986[4] && reverse_165986[3:0] == 4'h0, reverse_165986[3] && reverse_165986[2:0] == 3'h0, reverse_165986[2] && reverse_165986[1:0] == 2'h0, reverse_165986[1] && !reverse_165986[0], reverse_165986[0]};
  assign encode_165995 = {one_hot_165987[16] | one_hot_165987[17] | one_hot_165987[18] | one_hot_165987[19] | one_hot_165987[20] | one_hot_165987[21] | one_hot_165987[22] | one_hot_165987[23] | one_hot_165987[24] | one_hot_165987[25] | one_hot_165987[26] | one_hot_165987[27] | one_hot_165987[28], one_hot_165987[8] | one_hot_165987[9] | one_hot_165987[10] | one_hot_165987[11] | one_hot_165987[12] | one_hot_165987[13] | one_hot_165987[14] | one_hot_165987[15] | one_hot_165987[24] | one_hot_165987[25] | one_hot_165987[26] | one_hot_165987[27] | one_hot_165987[28], one_hot_165987[4] | one_hot_165987[5] | one_hot_165987[6] | one_hot_165987[7] | one_hot_165987[12] | one_hot_165987[13] | one_hot_165987[14] | one_hot_165987[15] | one_hot_165987[20] | one_hot_165987[21] | one_hot_165987[22] | one_hot_165987[23] | one_hot_165987[28], one_hot_165987[2] | one_hot_165987[3] | one_hot_165987[6] | one_hot_165987[7] | one_hot_165987[10] | one_hot_165987[11] | one_hot_165987[14] | one_hot_165987[15] | one_hot_165987[18] | one_hot_165987[19] | one_hot_165987[22] | one_hot_165987[23] | one_hot_165987[26] | one_hot_165987[27], one_hot_165987[1] | one_hot_165987[3] | one_hot_165987[5] | one_hot_165987[7] | one_hot_165987[9] | one_hot_165987[11] | one_hot_165987[13] | one_hot_165987[15] | one_hot_165987[17] | one_hot_165987[19] | one_hot_165987[21] | one_hot_165987[23] | one_hot_165987[25] | one_hot_165987[27]};
  assign encode_165996 = {one_hot_165988[16] | one_hot_165988[17] | one_hot_165988[18] | one_hot_165988[19] | one_hot_165988[20] | one_hot_165988[21] | one_hot_165988[22] | one_hot_165988[23] | one_hot_165988[24] | one_hot_165988[25] | one_hot_165988[26] | one_hot_165988[27] | one_hot_165988[28], one_hot_165988[8] | one_hot_165988[9] | one_hot_165988[10] | one_hot_165988[11] | one_hot_165988[12] | one_hot_165988[13] | one_hot_165988[14] | one_hot_165988[15] | one_hot_165988[24] | one_hot_165988[25] | one_hot_165988[26] | one_hot_165988[27] | one_hot_165988[28], one_hot_165988[4] | one_hot_165988[5] | one_hot_165988[6] | one_hot_165988[7] | one_hot_165988[12] | one_hot_165988[13] | one_hot_165988[14] | one_hot_165988[15] | one_hot_165988[20] | one_hot_165988[21] | one_hot_165988[22] | one_hot_165988[23] | one_hot_165988[28], one_hot_165988[2] | one_hot_165988[3] | one_hot_165988[6] | one_hot_165988[7] | one_hot_165988[10] | one_hot_165988[11] | one_hot_165988[14] | one_hot_165988[15] | one_hot_165988[18] | one_hot_165988[19] | one_hot_165988[22] | one_hot_165988[23] | one_hot_165988[26] | one_hot_165988[27], one_hot_165988[1] | one_hot_165988[3] | one_hot_165988[5] | one_hot_165988[7] | one_hot_165988[9] | one_hot_165988[11] | one_hot_165988[13] | one_hot_165988[15] | one_hot_165988[17] | one_hot_165988[19] | one_hot_165988[21] | one_hot_165988[23] | one_hot_165988[25] | one_hot_165988[27]};
  assign encode_165998 = {one_hot_165990[16] | one_hot_165990[17] | one_hot_165990[18] | one_hot_165990[19] | one_hot_165990[20] | one_hot_165990[21] | one_hot_165990[22] | one_hot_165990[23] | one_hot_165990[24] | one_hot_165990[25] | one_hot_165990[26] | one_hot_165990[27] | one_hot_165990[28], one_hot_165990[8] | one_hot_165990[9] | one_hot_165990[10] | one_hot_165990[11] | one_hot_165990[12] | one_hot_165990[13] | one_hot_165990[14] | one_hot_165990[15] | one_hot_165990[24] | one_hot_165990[25] | one_hot_165990[26] | one_hot_165990[27] | one_hot_165990[28], one_hot_165990[4] | one_hot_165990[5] | one_hot_165990[6] | one_hot_165990[7] | one_hot_165990[12] | one_hot_165990[13] | one_hot_165990[14] | one_hot_165990[15] | one_hot_165990[20] | one_hot_165990[21] | one_hot_165990[22] | one_hot_165990[23] | one_hot_165990[28], one_hot_165990[2] | one_hot_165990[3] | one_hot_165990[6] | one_hot_165990[7] | one_hot_165990[10] | one_hot_165990[11] | one_hot_165990[14] | one_hot_165990[15] | one_hot_165990[18] | one_hot_165990[19] | one_hot_165990[22] | one_hot_165990[23] | one_hot_165990[26] | one_hot_165990[27], one_hot_165990[1] | one_hot_165990[3] | one_hot_165990[5] | one_hot_165990[7] | one_hot_165990[9] | one_hot_165990[11] | one_hot_165990[13] | one_hot_165990[15] | one_hot_165990[17] | one_hot_165990[19] | one_hot_165990[21] | one_hot_165990[23] | one_hot_165990[25] | one_hot_165990[27]};
  assign encode_166000 = {one_hot_165992[16] | one_hot_165992[17] | one_hot_165992[18] | one_hot_165992[19] | one_hot_165992[20] | one_hot_165992[21] | one_hot_165992[22] | one_hot_165992[23] | one_hot_165992[24] | one_hot_165992[25] | one_hot_165992[26] | one_hot_165992[27] | one_hot_165992[28], one_hot_165992[8] | one_hot_165992[9] | one_hot_165992[10] | one_hot_165992[11] | one_hot_165992[12] | one_hot_165992[13] | one_hot_165992[14] | one_hot_165992[15] | one_hot_165992[24] | one_hot_165992[25] | one_hot_165992[26] | one_hot_165992[27] | one_hot_165992[28], one_hot_165992[4] | one_hot_165992[5] | one_hot_165992[6] | one_hot_165992[7] | one_hot_165992[12] | one_hot_165992[13] | one_hot_165992[14] | one_hot_165992[15] | one_hot_165992[20] | one_hot_165992[21] | one_hot_165992[22] | one_hot_165992[23] | one_hot_165992[28], one_hot_165992[2] | one_hot_165992[3] | one_hot_165992[6] | one_hot_165992[7] | one_hot_165992[10] | one_hot_165992[11] | one_hot_165992[14] | one_hot_165992[15] | one_hot_165992[18] | one_hot_165992[19] | one_hot_165992[22] | one_hot_165992[23] | one_hot_165992[26] | one_hot_165992[27], one_hot_165992[1] | one_hot_165992[3] | one_hot_165992[5] | one_hot_165992[7] | one_hot_165992[9] | one_hot_165992[11] | one_hot_165992[13] | one_hot_165992[15] | one_hot_165992[17] | one_hot_165992[19] | one_hot_165992[21] | one_hot_165992[23] | one_hot_165992[25] | one_hot_165992[27]};
  assign encode_166002 = {one_hot_165994[16] | one_hot_165994[17] | one_hot_165994[18] | one_hot_165994[19] | one_hot_165994[20] | one_hot_165994[21] | one_hot_165994[22] | one_hot_165994[23] | one_hot_165994[24] | one_hot_165994[25] | one_hot_165994[26] | one_hot_165994[27] | one_hot_165994[28], one_hot_165994[8] | one_hot_165994[9] | one_hot_165994[10] | one_hot_165994[11] | one_hot_165994[12] | one_hot_165994[13] | one_hot_165994[14] | one_hot_165994[15] | one_hot_165994[24] | one_hot_165994[25] | one_hot_165994[26] | one_hot_165994[27] | one_hot_165994[28], one_hot_165994[4] | one_hot_165994[5] | one_hot_165994[6] | one_hot_165994[7] | one_hot_165994[12] | one_hot_165994[13] | one_hot_165994[14] | one_hot_165994[15] | one_hot_165994[20] | one_hot_165994[21] | one_hot_165994[22] | one_hot_165994[23] | one_hot_165994[28], one_hot_165994[2] | one_hot_165994[3] | one_hot_165994[6] | one_hot_165994[7] | one_hot_165994[10] | one_hot_165994[11] | one_hot_165994[14] | one_hot_165994[15] | one_hot_165994[18] | one_hot_165994[19] | one_hot_165994[22] | one_hot_165994[23] | one_hot_165994[26] | one_hot_165994[27], one_hot_165994[1] | one_hot_165994[3] | one_hot_165994[5] | one_hot_165994[7] | one_hot_165994[9] | one_hot_165994[11] | one_hot_165994[13] | one_hot_165994[15] | one_hot_165994[17] | one_hot_165994[19] | one_hot_165994[21] | one_hot_165994[23] | one_hot_165994[25] | one_hot_165994[27]};
  assign cancel__15 = |encode_165989[4:1];
  assign carry_bit__14 = xbs_fraction__14[27];
  assign result_fraction__508 = 23'h00_0000;
  assign cancel__30 = |encode_165991[4:1];
  assign carry_bit__30 = xbs_fraction__29[27];
  assign result_fraction__575 = 23'h00_0000;
  assign cancel__49 = |encode_165993[4:1];
  assign carry_bit__49 = xbs_fraction__47[27];
  assign result_fraction__640 = 23'h00_0000;
  assign cancel__68 = |encode_165995[4:1];
  assign carry_bit__68 = xbs_fraction__65[27];
  assign result_fraction__715 = 23'h00_0000;
  assign cancel__6 = |encode_165996[4:1];
  assign carry_bit__6 = xbs_fraction__6[27];
  assign result_fraction__509 = 23'h00_0000;
  assign leading_zeroes__14 = {result_fraction__508, encode_165989};
  assign cancel__31 = |encode_165998[4:1];
  assign carry_bit__31 = xbs_fraction__30[27];
  assign result_fraction__576 = 23'h00_0000;
  assign leading_zeroes__30 = {result_fraction__575, encode_165991};
  assign cancel__50 = |encode_166000[4:1];
  assign carry_bit__50 = xbs_fraction__48[27];
  assign result_fraction__641 = 23'h00_0000;
  assign leading_zeroes__49 = {result_fraction__640, encode_165993};
  assign cancel__69 = |encode_166002[4:1];
  assign carry_bit__69 = xbs_fraction__66[27];
  assign result_fraction__716 = 23'h00_0000;
  assign leading_zeroes__68 = {result_fraction__715, encode_165995};
  assign leading_zeroes__6 = {result_fraction__509, encode_165996};
  assign carry_fraction__28 = xbs_fraction__14[27:1];
  assign add_166070 = leading_zeroes__14 + 28'hfff_ffff;
  assign leading_zeroes__31 = {result_fraction__576, encode_165998};
  assign carry_fraction__59 = xbs_fraction__29[27:1];
  assign add_166083 = leading_zeroes__30 + 28'hfff_ffff;
  assign leading_zeroes__50 = {result_fraction__641, encode_166000};
  assign carry_fraction__97 = xbs_fraction__47[27:1];
  assign add_166096 = leading_zeroes__49 + 28'hfff_ffff;
  assign array_index_166097 = in_img_unflattened[4'hc];
  assign leading_zeroes__69 = {result_fraction__716, encode_166002};
  assign carry_fraction__135 = xbs_fraction__65[27:1];
  assign add_166110 = leading_zeroes__68 + 28'hfff_ffff;
  assign array_index_166111 = in_img_unflattened[4'hd];
  assign carry_fraction__11 = xbs_fraction__6[27:1];
  assign add_166118 = leading_zeroes__6 + 28'hfff_ffff;
  assign concat_166119 = {~(carry_bit__14 | cancel__15), ~(carry_bit__14 | ~cancel__15), ~(~carry_bit__14 | cancel__15)};
  assign carry_fraction__29 = carry_fraction__28 | {26'h000_0000, xbs_fraction__14[0]};
  assign cancel_fraction__14 = add_166070 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__14[26:0] << add_166070;
  assign result_sign__599 = 1'h0;
  assign carry_fraction__60 = xbs_fraction__30[27:1];
  assign add_166129 = leading_zeroes__31 + 28'hfff_ffff;
  assign concat_166130 = {~(carry_bit__30 | cancel__30), ~(carry_bit__30 | ~cancel__30), ~(~carry_bit__30 | cancel__30)};
  assign carry_fraction__61 = carry_fraction__59 | {26'h000_0000, xbs_fraction__29[0]};
  assign cancel_fraction__30 = add_166083 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__29[26:0] << add_166083;
  assign result_sign__705 = 1'h0;
  assign carry_fraction__98 = xbs_fraction__48[27:1];
  assign add_166140 = leading_zeroes__50 + 28'hfff_ffff;
  assign concat_166141 = {~(carry_bit__49 | cancel__49), ~(carry_bit__49 | ~cancel__49), ~(~carry_bit__49 | cancel__49)};
  assign carry_fraction__99 = carry_fraction__97 | {26'h000_0000, xbs_fraction__47[0]};
  assign cancel_fraction__49 = add_166096 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__47[26:0] << add_166096;
  assign result_sign__630 = 1'h0;
  assign x_bexp__381 = array_index_166097[30:23];
  assign carry_fraction__136 = xbs_fraction__66[27:1];
  assign add_166152 = leading_zeroes__69 + 28'hfff_ffff;
  assign concat_166153 = {~(carry_bit__68 | cancel__68), ~(carry_bit__68 | ~cancel__68), ~(~carry_bit__68 | cancel__68)};
  assign carry_fraction__137 = carry_fraction__135 | {26'h000_0000, xbs_fraction__65[0]};
  assign cancel_fraction__68 = add_166110 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__65[26:0] << add_166110;
  assign result_sign__738 = 1'h0;
  assign x_bexp__525 = array_index_166111[30:23];
  assign concat_166158 = {~(carry_bit__6 | cancel__6), ~(carry_bit__6 | ~cancel__6), ~(~carry_bit__6 | cancel__6)};
  assign carry_fraction__12 = carry_fraction__11 | {26'h000_0000, xbs_fraction__6[0]};
  assign cancel_fraction__6 = add_166118 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__6[26:0] << add_166118;
  assign shifted_fraction__14 = carry_fraction__29 & {27{concat_166119[0]}} | cancel_fraction__14 & {27{concat_166119[1]}} | xbs_fraction__14[26:0] & {27{concat_166119[2]}};
  assign concat_166164 = {~(carry_bit__31 | cancel__31), ~(carry_bit__31 | ~cancel__31), ~(~carry_bit__31 | cancel__31)};
  assign carry_fraction__62 = carry_fraction__60 | {26'h000_0000, xbs_fraction__30[0]};
  assign cancel_fraction__31 = add_166129 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__30[26:0] << add_166129;
  assign shifted_fraction__30 = carry_fraction__61 & {27{concat_166130[0]}} | cancel_fraction__30 & {27{concat_166130[1]}} | xbs_fraction__29[26:0] & {27{concat_166130[2]}};
  assign concat_166170 = {~(carry_bit__50 | cancel__50), ~(carry_bit__50 | ~cancel__50), ~(~carry_bit__50 | cancel__50)};
  assign carry_fraction__100 = carry_fraction__98 | {26'h000_0000, xbs_fraction__48[0]};
  assign cancel_fraction__50 = add_166140 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__48[26:0] << add_166140;
  assign shifted_fraction__49 = carry_fraction__99 & {27{concat_166141[0]}} | cancel_fraction__49 & {27{concat_166141[1]}} | xbs_fraction__47[26:0] & {27{concat_166141[2]}};
  assign concat_166176 = {~(carry_bit__69 | cancel__69), ~(carry_bit__69 | ~cancel__69), ~(~carry_bit__69 | cancel__69)};
  assign carry_fraction__138 = carry_fraction__136 | {26'h000_0000, xbs_fraction__66[0]};
  assign cancel_fraction__69 = add_166152 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__66[26:0] << add_166152;
  assign shifted_fraction__68 = carry_fraction__137 & {27{concat_166153[0]}} | cancel_fraction__68 & {27{concat_166153[1]}} | xbs_fraction__65[26:0] & {27{concat_166153[2]}};
  assign shifted_fraction__6 = carry_fraction__12 & {27{concat_166158[0]}} | cancel_fraction__6 & {27{concat_166158[1]}} | xbs_fraction__6[26:0] & {27{concat_166158[2]}};
  assign result_sign__1042 = 1'h0;
  assign result_sign__435 = 1'h0;
  assign add_166186 = {result_sign__599, x_bexp__334} + 9'h07f;
  assign shifted_fraction__31 = carry_fraction__62 & {27{concat_166164[0]}} | cancel_fraction__31 & {27{concat_166164[1]}} | xbs_fraction__30[26:0] & {27{concat_166164[2]}};
  assign result_sign__1043 = 1'h0;
  assign result_sign__532 = 1'h0;
  assign add_166191 = {result_sign__705, x_bexp__478} + 9'h07f;
  assign shifted_fraction__50 = carry_fraction__100 & {27{concat_166170[0]}} | cancel_fraction__50 & {27{concat_166170[1]}} | xbs_fraction__48[26:0] & {27{concat_166170[2]}};
  assign result_sign__1044 = 1'h0;
  assign result_sign__632 = 1'h0;
  assign add_166196 = {result_sign__630, x_bexp__381} + 9'h07f;
  assign x_bexp__760 = 8'h00;
  assign result_sign__628 = 1'h0;
  assign x_fraction__381 = array_index_166097[22:0];
  assign shifted_fraction__69 = carry_fraction__138 & {27{concat_166176[0]}} | cancel_fraction__69 & {27{concat_166176[1]}} | xbs_fraction__66[26:0] & {27{concat_166176[2]}};
  assign result_sign__1045 = 1'h0;
  assign result_sign__740 = 1'h0;
  assign add_166204 = {result_sign__738, x_bexp__525} + 9'h07f;
  assign x_bexp__761 = 8'h00;
  assign result_sign__736 = 1'h0;
  assign x_fraction__525 = array_index_166111[22:0];
  assign result_sign__1046 = 1'h0;
  assign normal_chunk__14 = shifted_fraction__14[2:0];
  assign fraction_shift__245 = 3'h4;
  assign half_way_chunk__14 = shifted_fraction__14[3:2];
  assign result_sign__1047 = 1'h0;
  assign normal_chunk__30 = shifted_fraction__30[2:0];
  assign fraction_shift__280 = 3'h4;
  assign half_way_chunk__30 = shifted_fraction__30[3:2];
  assign result_sign__1048 = 1'h0;
  assign normal_chunk__49 = shifted_fraction__49[2:0];
  assign fraction_shift__315 = 3'h4;
  assign half_way_chunk__49 = shifted_fraction__49[3:2];
  assign ne_166238 = x_bexp__381 != x_bexp__760;
  assign result_sign__1049 = 1'h0;
  assign normal_chunk__68 = shifted_fraction__68[2:0];
  assign fraction_shift__350 = 3'h4;
  assign half_way_chunk__68 = shifted_fraction__68[3:2];
  assign ne_166251 = x_bexp__525 != x_bexp__761;
  assign normal_chunk__6 = shifted_fraction__6[2:0];
  assign fraction_shift__246 = 3'h4;
  assign half_way_chunk__6 = shifted_fraction__6[3:2];
  assign result_sign__432 = 1'h0;
  assign add_166263 = {result_sign__1042, shifted_fraction__14[26:3]} + 25'h000_0001;
  assign exp__60 = {result_sign__435, add_166186} + 10'h381;
  assign normal_chunk__31 = shifted_fraction__31[2:0];
  assign fraction_shift__281 = 3'h4;
  assign half_way_chunk__31 = shifted_fraction__31[3:2];
  assign result_sign__529 = 1'h0;
  assign add_166274 = {result_sign__1043, shifted_fraction__30[26:3]} + 25'h000_0001;
  assign exp__131 = {result_sign__532, add_166191} + 10'h381;
  assign normal_chunk__50 = shifted_fraction__50[2:0];
  assign fraction_shift__316 = 3'h4;
  assign half_way_chunk__50 = shifted_fraction__50[3:2];
  assign result_sign__627 = 1'h0;
  assign add_166285 = {result_sign__1044, shifted_fraction__49[26:3]} + 25'h000_0001;
  assign exp__213 = {result_sign__632, add_166196} + 10'h381;
  assign x_fraction__383 = {result_sign__628, x_fraction__381} | 24'h80_0000;
  assign normal_chunk__69 = shifted_fraction__69[2:0];
  assign fraction_shift__351 = 3'h4;
  assign half_way_chunk__69 = shifted_fraction__69[3:2];
  assign result_sign__735 = 1'h0;
  assign add_166299 = {result_sign__1045, shifted_fraction__68[26:3]} + 25'h000_0001;
  assign exp__295 = {result_sign__740, add_166204} + 10'h381;
  assign sign_ext_166301 = {10{ne_166251}};
  assign x_fraction__527 = {result_sign__736, x_fraction__525} | 24'h80_0000;
  assign result_sign__433 = 1'h0;
  assign add_166307 = {result_sign__1046, shifted_fraction__6[26:3]} + 25'h000_0001;
  assign do_round_up__29 = normal_chunk__14 > fraction_shift__245 | half_way_chunk__14 == 2'h3;
  assign exp__61 = exp__60 & sign_ext_161429;
  assign result_sign__530 = 1'h0;
  assign add_166316 = {result_sign__1047, shifted_fraction__31[26:3]} + 25'h000_0001;
  assign do_round_up__62 = normal_chunk__30 > fraction_shift__280 | half_way_chunk__30 == 2'h3;
  assign exp__133 = exp__131 & sign_ext_161440;
  assign result_sign__629 = 1'h0;
  assign add_166325 = {result_sign__1048, shifted_fraction__50[26:3]} + 25'h000_0001;
  assign do_round_up__101 = normal_chunk__49 > fraction_shift__315 | half_way_chunk__49 == 2'h3;
  assign exp__215 = exp__213 & {10{ne_166238}};
  assign x_fraction__385 = x_fraction__383 & {24{ne_166238}};
  assign result_sign__820 = 1'h0;
  assign result_sign__821 = 1'h0;
  assign result_sign__737 = 1'h0;
  assign add_166337 = {result_sign__1049, shifted_fraction__69[26:3]} + 25'h000_0001;
  assign do_round_up__140 = normal_chunk__68 > fraction_shift__350 | half_way_chunk__68 == 2'h3;
  assign exp__297 = exp__295 & sign_ext_166301;
  assign x_fraction__529 = x_fraction__527 & {24{ne_166251}};
  assign result_sign__822 = 1'h0;
  assign result_sign__823 = 1'h0;
  assign do_round_up__12 = normal_chunk__6 > fraction_shift__246 | half_way_chunk__6 == 2'h3;
  assign rounded_fraction__14 = do_round_up__29 ? {add_166263, normal_chunk__14} : {result_sign__432, shifted_fraction__14};
  assign do_round_up__63 = normal_chunk__31 > fraction_shift__281 | half_way_chunk__31 == 2'h3;
  assign rounded_fraction__30 = do_round_up__62 ? {add_166274, normal_chunk__30} : {result_sign__529, shifted_fraction__30};
  assign do_round_up__102 = normal_chunk__50 > fraction_shift__316 | half_way_chunk__50 == 2'h3;
  assign rounded_fraction__49 = do_round_up__101 ? {add_166285, normal_chunk__49} : {result_sign__627, shifted_fraction__49};
  assign do_round_up__141 = normal_chunk__69 > fraction_shift__351 | half_way_chunk__69 == 2'h3;
  assign rounded_fraction__68 = do_round_up__140 ? {add_166299, normal_chunk__68} : {result_sign__735, shifted_fraction__68};
  assign concat_166368 = {x_fraction__529, result_sign__822};
  assign concat_166369 = {result_sign__823, x_fraction__529};
  assign rounded_fraction__6 = do_round_up__12 ? {add_166307, normal_chunk__6} : {result_sign__433, shifted_fraction__6};
  assign result_sign__434 = 1'h0;
  assign x_bexp__584 = 8'h00;
  assign rounding_carry__14 = rounded_fraction__14[27];
  assign sel_166374 = $signed(exp__61) <= $signed(10'h000) ? concat_161486 : concat_161485;
  assign rounded_fraction__31 = do_round_up__63 ? {add_166316, normal_chunk__31} : {result_sign__530, shifted_fraction__31};
  assign result_sign__531 = 1'h0;
  assign x_bexp__602 = 8'h00;
  assign rounding_carry__30 = rounded_fraction__30[27];
  assign sel_166379 = $signed(exp__133) <= $signed(10'h000) ? concat_161493 : concat_161492;
  assign rounded_fraction__50 = do_round_up__102 ? {add_166325, normal_chunk__50} : {result_sign__629, shifted_fraction__50};
  assign result_sign__631 = 1'h0;
  assign x_bexp__620 = 8'h00;
  assign rounding_carry__49 = rounded_fraction__49[27];
  assign sel_166384 = $signed(exp__215) <= $signed(10'h000) ? {result_sign__821, x_fraction__385} : {x_fraction__385, result_sign__820};
  assign rounded_fraction__69 = do_round_up__141 ? {add_166337, normal_chunk__69} : {result_sign__737, shifted_fraction__69};
  assign result_sign__739 = 1'h0;
  assign x_bexp__638 = 8'h00;
  assign rounding_carry__68 = rounded_fraction__68[27];
  assign sel_166389 = $signed(exp__297) <= $signed(10'h000) ? concat_166369 : concat_166368;
  assign result_sign__436 = 1'h0;
  assign x_bexp__585 = 8'h00;
  assign rounding_carry__6 = rounded_fraction__6[27];
  assign result_sign__932 = 1'h0;
  assign fraction__140 = sel_166374[23:1];
  assign result_sign__533 = 1'h0;
  assign x_bexp__603 = 8'h00;
  assign rounding_carry__31 = rounded_fraction__31[27];
  assign result_sign__938 = 1'h0;
  assign fraction__298 = sel_166379[23:1];
  assign result_sign__633 = 1'h0;
  assign x_bexp__621 = 8'h00;
  assign rounding_carry__50 = rounded_fraction__50[27];
  assign result_sign__945 = 1'h0;
  assign fraction__477 = sel_166384[23:1];
  assign result_sign__741 = 1'h0;
  assign x_bexp__639 = 8'h00;
  assign rounding_carry__69 = rounded_fraction__69[27];
  assign result_sign__953 = 1'h0;
  assign fraction__656 = sel_166389[23:1];
  assign result_sign__437 = 1'h0;
  assign add_166421 = {result_sign__434, x_bexp__118} + {x_bexp__584, rounding_carry__14};
  assign fraction__141 = {result_sign__932, fraction__140};
  assign result_sign__534 = 1'h0;
  assign add_166431 = {result_sign__531, x_bexp__235} + {x_bexp__602, rounding_carry__30};
  assign fraction__300 = {result_sign__938, fraction__298};
  assign result_sign__634 = 1'h0;
  assign add_166441 = {result_sign__631, x_bexp__379} + {x_bexp__620, rounding_carry__49};
  assign fraction__479 = {result_sign__945, fraction__477};
  assign result_sign__742 = 1'h0;
  assign add_166451 = {result_sign__739, x_bexp__523} + {x_bexp__638, rounding_carry__68};
  assign fraction__658 = {result_sign__953, fraction__656};
  assign result_sign__438 = 1'h0;
  assign add_166459 = {result_sign__436, x_bexp__46} + {x_bexp__585, rounding_carry__6};
  assign do_round_up__30 = sel_166374[0] & sel_166374[1];
  assign add_166468 = fraction__141 + 24'h00_0001;
  assign result_sign__535 = 1'h0;
  assign add_166470 = {result_sign__533, x_bexp__236} + {x_bexp__603, rounding_carry__31};
  assign do_round_up__64 = sel_166379[0] & sel_166379[1];
  assign add_166479 = fraction__300 + 24'h00_0001;
  assign result_sign__635 = 1'h0;
  assign add_166481 = {result_sign__633, x_bexp__380} + {x_bexp__621, rounding_carry__50};
  assign do_round_up__103 = sel_166384[0] & sel_166384[1];
  assign add_166490 = fraction__479 + 24'h00_0001;
  assign result_sign__743 = 1'h0;
  assign add_166492 = {result_sign__741, x_bexp__524} + {x_bexp__639, rounding_carry__69};
  assign do_round_up__142 = sel_166389[0] & sel_166389[1];
  assign add_166501 = fraction__658 + 24'h00_0001;
  assign add_166507 = {result_sign__437, add_166421} + 10'h001;
  assign fraction__142 = do_round_up__30 ? add_166468 : fraction__141;
  assign add_166517 = {result_sign__534, add_166431} + 10'h001;
  assign fraction__302 = do_round_up__64 ? add_166479 : fraction__300;
  assign add_166527 = {result_sign__634, add_166441} + 10'h001;
  assign fraction__481 = do_round_up__103 ? add_166490 : fraction__479;
  assign add_166537 = {result_sign__742, add_166451} + 10'h001;
  assign fraction__660 = do_round_up__142 ? add_166501 : fraction__658;
  assign add_166542 = {result_sign__438, add_166459} + 10'h001;
  assign wide_exponent__42 = add_166507 - {5'h00, encode_165989};
  assign add_166548 = exp__61 + 10'h001;
  assign add_166549 = {result_sign__535, add_166470} + 10'h001;
  assign wide_exponent__88 = add_166517 - {5'h00, encode_165991};
  assign add_166555 = exp__133 + 10'h001;
  assign add_166556 = {result_sign__635, add_166481} + 10'h001;
  assign wide_exponent__145 = add_166527 - {5'h00, encode_165993};
  assign add_166562 = exp__215 + 10'h001;
  assign add_166563 = {result_sign__743, add_166492} + 10'h001;
  assign wide_exponent__202 = add_166537 - {5'h00, encode_165995};
  assign add_166569 = exp__297 + 10'h001;
  assign wide_exponent__16 = add_166542 - {5'h00, encode_165996};
  assign wide_exponent__43 = wide_exponent__42 & {10{add_165914 != 26'h000_0000 | xddend_y__14[2:0] != 3'h0}};
  assign exp__63 = fraction__142[23] ? add_166548 : exp__61;
  assign wide_exponent__89 = add_166549 - {5'h00, encode_165998};
  assign wide_exponent__90 = wide_exponent__88 & {10{add_165917 != 26'h000_0000 | xddend_y__29[2:0] != 3'h0}};
  assign exp__137 = fraction__302[23] ? add_166555 : exp__133;
  assign wide_exponent__146 = add_166556 - {5'h00, encode_166000};
  assign wide_exponent__147 = wide_exponent__145 & {10{add_165920 != 26'h000_0000 | xddend_y__47[2:0] != 3'h0}};
  assign exp__219 = fraction__481[23] ? add_166562 : exp__215;
  assign wide_exponent__203 = add_166563 - {5'h00, encode_166002};
  assign wide_exponent__204 = wide_exponent__202 & {10{add_165923 != 26'h000_0000 | xddend_y__65[2:0] != 3'h0}};
  assign exp__301 = fraction__660[23] ? add_166569 : exp__297;
  assign wide_exponent__17 = wide_exponent__16 & {10{add_165924 != 26'h000_0000 | xddend_y__6[2:0] != 3'h0}};
  assign high_exp__373 = 8'hff;
  assign result_fraction__779 = 23'h00_0000;
  assign high_exp__374 = 8'hff;
  assign result_fraction__780 = 23'h00_0000;
  assign high_exp__110 = 8'hff;
  assign result_fraction__510 = 23'h00_0000;
  assign high_exp__111 = 8'hff;
  assign result_fraction__511 = 23'h00_0000;
  assign wide_exponent__91 = wide_exponent__89 & {10{add_165927 != 26'h000_0000 | xddend_y__30[2:0] != 3'h0}};
  assign high_exp__405 = 8'hff;
  assign result_fraction__812 = 23'h00_0000;
  assign high_exp__406 = 8'hff;
  assign result_fraction__813 = 23'h00_0000;
  assign high_exp__175 = 8'hff;
  assign result_fraction__577 = 23'h00_0000;
  assign high_exp__176 = 8'hff;
  assign result_fraction__578 = 23'h00_0000;
  assign wide_exponent__148 = wide_exponent__146 & {10{add_165930 != 26'h000_0000 | xddend_y__48[2:0] != 3'h0}};
  assign high_exp__437 = 8'hff;
  assign result_fraction__845 = 23'h00_0000;
  assign high_exp__438 = 8'hff;
  assign result_fraction__846 = 23'h00_0000;
  assign high_exp__241 = 8'hff;
  assign result_fraction__642 = 23'h00_0000;
  assign high_exp__242 = 8'hff;
  assign result_fraction__643 = 23'h00_0000;
  assign wide_exponent__205 = wide_exponent__203 & {10{add_165933 != 26'h000_0000 | xddend_y__66[2:0] != 3'h0}};
  assign high_exp__469 = 8'hff;
  assign result_fraction__878 = 23'h00_0000;
  assign high_exp__470 = 8'hff;
  assign result_fraction__879 = 23'h00_0000;
  assign high_exp__313 = 8'hff;
  assign result_fraction__717 = 23'h00_0000;
  assign high_exp__314 = 8'hff;
  assign result_fraction__718 = 23'h00_0000;
  assign high_exp__359 = 8'hff;
  assign result_fraction__764 = 23'h00_0000;
  assign high_exp__360 = 8'hff;
  assign result_fraction__765 = 23'h00_0000;
  assign high_exp__112 = 8'hff;
  assign result_fraction__512 = 23'h00_0000;
  assign high_exp__113 = 8'hff;
  assign result_fraction__513 = 23'h00_0000;
  assign ne_166645 = x_fraction__118 != result_fraction__779;
  assign ne_166647 = prod_fraction__42 != result_fraction__780;
  assign eq_166648 = x_bexp__118 == high_exp__110;
  assign eq_166649 = x_fraction__118 == result_fraction__510;
  assign eq_166650 = prod_bexp__58 == high_exp__111;
  assign eq_166651 = prod_fraction__42 == result_fraction__511;
  assign result_exp__45 = exp__63[8:0];
  assign high_exp__391 = 8'hff;
  assign result_fraction__797 = 23'h00_0000;
  assign high_exp__392 = 8'hff;
  assign result_fraction__798 = 23'h00_0000;
  assign high_exp__177 = 8'hff;
  assign result_fraction__579 = 23'h00_0000;
  assign high_exp__178 = 8'hff;
  assign result_fraction__580 = 23'h00_0000;
  assign ne_166665 = x_fraction__235 != result_fraction__812;
  assign ne_166667 = prod_fraction__85 != result_fraction__813;
  assign eq_166668 = x_bexp__235 == high_exp__175;
  assign eq_166669 = x_fraction__235 == result_fraction__577;
  assign eq_166670 = prod_bexp__115 == high_exp__176;
  assign eq_166671 = prod_fraction__85 == result_fraction__578;
  assign result_exp__97 = exp__137[8:0];
  assign high_exp__423 = 8'hff;
  assign result_fraction__830 = 23'h00_0000;
  assign high_exp__424 = 8'hff;
  assign result_fraction__831 = 23'h00_0000;
  assign high_exp__243 = 8'hff;
  assign result_fraction__644 = 23'h00_0000;
  assign high_exp__244 = 8'hff;
  assign result_fraction__645 = 23'h00_0000;
  assign ne_166685 = x_fraction__379 != result_fraction__845;
  assign ne_166687 = prod_fraction__139 != result_fraction__846;
  assign eq_166688 = x_bexp__379 == high_exp__241;
  assign eq_166689 = x_fraction__379 == result_fraction__642;
  assign eq_166690 = prod_bexp__187 == high_exp__242;
  assign eq_166691 = prod_fraction__139 == result_fraction__643;
  assign result_exp__157 = exp__219[8:0];
  assign high_exp__455 = 8'hff;
  assign result_fraction__863 = 23'h00_0000;
  assign high_exp__456 = 8'hff;
  assign result_fraction__864 = 23'h00_0000;
  assign high_exp__315 = 8'hff;
  assign result_fraction__719 = 23'h00_0000;
  assign high_exp__316 = 8'hff;
  assign result_fraction__720 = 23'h00_0000;
  assign ne_166705 = x_fraction__523 != result_fraction__878;
  assign ne_166707 = prod_fraction__193 != result_fraction__879;
  assign eq_166708 = x_bexp__523 == high_exp__313;
  assign eq_166709 = x_fraction__523 == result_fraction__717;
  assign eq_166710 = prod_bexp__259 == high_exp__314;
  assign eq_166711 = prod_fraction__193 == result_fraction__718;
  assign result_exp__217 = exp__301[8:0];
  assign ne_166716 = x_fraction__46 != result_fraction__764;
  assign ne_166718 = prod_fraction__16 != result_fraction__765;
  assign eq_166719 = x_bexp__46 == high_exp__112;
  assign eq_166720 = x_fraction__46 == result_fraction__512;
  assign eq_166721 = prod_bexp__22 == high_exp__113;
  assign eq_166722 = prod_fraction__16 == result_fraction__513;
  assign result_exp__46 = result_exp__45 & {9{$signed(exp__63) > $signed(10'h000)}};
  assign ne_166732 = x_fraction__236 != result_fraction__797;
  assign ne_166734 = prod_fraction__86 != result_fraction__798;
  assign eq_166735 = x_bexp__236 == high_exp__177;
  assign eq_166736 = x_fraction__236 == result_fraction__579;
  assign eq_166737 = prod_bexp__116 == high_exp__178;
  assign eq_166738 = prod_fraction__86 == result_fraction__580;
  assign result_exp__99 = result_exp__97 & {9{$signed(exp__137) > $signed(10'h000)}};
  assign ne_166748 = x_fraction__380 != result_fraction__830;
  assign ne_166750 = prod_fraction__140 != result_fraction__831;
  assign eq_166751 = x_bexp__380 == high_exp__243;
  assign eq_166752 = x_fraction__380 == result_fraction__644;
  assign eq_166753 = prod_bexp__188 == high_exp__244;
  assign eq_166754 = prod_fraction__140 == result_fraction__645;
  assign high_exp__247 = 8'hff;
  assign result_fraction__647 = 23'h00_0000;
  assign result_fraction__646 = 23'h00_0000;
  assign result_exp__159 = result_exp__157 & {9{$signed(exp__219) > $signed(10'h000)}};
  assign ne_166767 = x_fraction__524 != result_fraction__863;
  assign ne_166769 = prod_fraction__194 != result_fraction__864;
  assign eq_166770 = x_bexp__524 == high_exp__315;
  assign eq_166771 = x_fraction__524 == result_fraction__719;
  assign eq_166772 = prod_bexp__260 == high_exp__316;
  assign eq_166773 = prod_fraction__194 == result_fraction__720;
  assign high_exp__319 = 8'hff;
  assign result_fraction__722 = 23'h00_0000;
  assign result_fraction__721 = 23'h00_0000;
  assign result_exp__219 = result_exp__217 & {9{$signed(exp__301) > $signed(10'h000)}};
  assign wide_exponent__44 = wide_exponent__43[8:0] & {9{~wide_exponent__43[9]}};
  assign has_pos_inf__14 = ~(x_bexp__118 != high_exp__373 | ne_166645 | x_sign__30) | ~(prod_bexp__58 != high_exp__374 | ne_166647 | prod_sign__14);
  assign has_neg_inf__14 = eq_166648 & eq_166649 & x_sign__30 | eq_166650 & eq_166651 & prod_sign__14;
  assign wide_exponent__92 = wide_exponent__90[8:0] & {9{~wide_exponent__90[9]}};
  assign has_pos_inf__30 = ~(x_bexp__235 != high_exp__405 | ne_166665 | x_sign__59) | ~(prod_bexp__115 != high_exp__406 | ne_166667 | prod_sign__29);
  assign has_neg_inf__30 = eq_166668 & eq_166669 & x_sign__59 | eq_166670 & eq_166671 & prod_sign__29;
  assign wide_exponent__149 = wide_exponent__147[8:0] & {9{~wide_exponent__147[9]}};
  assign has_pos_inf__49 = ~(x_bexp__379 != high_exp__437 | ne_166685 | x_sign__95) | ~(prod_bexp__187 != high_exp__438 | ne_166687 | prod_sign__47);
  assign has_neg_inf__49 = eq_166688 & eq_166689 & x_sign__95 | eq_166690 & eq_166691 & prod_sign__47;
  assign eq_166813 = x_bexp__381 == high_exp__247;
  assign ne_166814 = x_fraction__381 != result_fraction__647;
  assign wide_exponent__206 = wide_exponent__204[8:0] & {9{~wide_exponent__204[9]}};
  assign has_pos_inf__68 = ~(x_bexp__523 != high_exp__469 | ne_166705 | x_sign__131) | ~(prod_bexp__259 != high_exp__470 | ne_166707 | prod_sign__65);
  assign has_neg_inf__68 = eq_166708 & eq_166709 & x_sign__131 | eq_166710 & eq_166711 & prod_sign__65;
  assign is_result_nan__108 = x_bexp__525 == high_exp__319;
  assign ne_166827 = x_fraction__525 != result_fraction__722;
  assign wide_exponent__18 = wide_exponent__17[8:0] & {9{~wide_exponent__17[9]}};
  assign has_pos_inf__6 = ~(x_bexp__46 != high_exp__359 | ne_166716 | x_sign__12) | ~(prod_bexp__22 != high_exp__360 | ne_166718 | prod_sign__6);
  assign has_neg_inf__6 = eq_166719 & eq_166720 & x_sign__12 | eq_166721 & eq_166722 & prod_sign__6;
  assign and_reduce_166841 = &result_exp__46[7:0];
  assign wide_exponent__93 = wide_exponent__91[8:0] & {9{~wide_exponent__91[9]}};
  assign has_pos_inf__31 = ~(x_bexp__236 != high_exp__391 | ne_166732 | x_sign__60) | ~(prod_bexp__116 != high_exp__392 | ne_166734 | prod_sign__30);
  assign has_neg_inf__31 = eq_166735 & eq_166736 & x_sign__60 | eq_166737 & eq_166738 & prod_sign__30;
  assign and_reduce_166853 = &result_exp__99[7:0];
  assign wide_exponent__150 = wide_exponent__148[8:0] & {9{~wide_exponent__148[9]}};
  assign has_pos_inf__50 = ~(x_bexp__380 != high_exp__423 | ne_166748 | x_sign__96) | ~(prod_bexp__188 != high_exp__424 | ne_166750 | prod_sign__48);
  assign has_neg_inf__50 = eq_166751 & eq_166752 & x_sign__96 | eq_166753 & eq_166754 & prod_sign__48;
  assign is_result_nan__103 = eq_166813 & ne_166814;
  assign has_inf_arg__53 = eq_166813 & x_fraction__381 == result_fraction__646;
  assign and_reduce_166867 = &result_exp__159[7:0];
  assign wide_exponent__207 = wide_exponent__205[8:0] & {9{~wide_exponent__205[9]}};
  assign has_pos_inf__69 = ~(x_bexp__524 != high_exp__455 | ne_166767 | x_sign__132) | ~(prod_bexp__260 != high_exp__456 | ne_166769 | prod_sign__66);
  assign has_neg_inf__69 = eq_166770 & eq_166771 & x_sign__132 | eq_166772 & eq_166773 & prod_sign__66;
  assign is_result_nan__142 = is_result_nan__108 & ne_166827;
  assign has_inf_arg__73 = is_result_nan__108 & x_fraction__525 == result_fraction__721;
  assign and_reduce_166881 = &result_exp__219[7:0];
  assign is_result_nan__29 = eq_166648 & ne_166645 | eq_166650 & ne_166647 | has_pos_inf__14 & has_neg_inf__14;
  assign is_operand_inf__14 = eq_166648 & eq_166649 | eq_166650 & eq_166651;
  assign and_reduce_166895 = &wide_exponent__44[7:0];
  assign high_exp__116 = 8'hff;
  assign is_result_nan__62 = eq_166668 & ne_166665 | eq_166670 & ne_166667 | has_pos_inf__30 & has_neg_inf__30;
  assign is_operand_inf__30 = eq_166668 & eq_166669 | eq_166670 & eq_166671;
  assign and_reduce_166911 = &wide_exponent__92[7:0];
  assign high_exp__181 = 8'hff;
  assign is_result_nan__101 = eq_166688 & ne_166685 | eq_166690 & ne_166687 | has_pos_inf__49 & has_neg_inf__49;
  assign is_operand_inf__49 = eq_166688 & eq_166689 | eq_166690 & eq_166691;
  assign and_reduce_166927 = &wide_exponent__149[7:0];
  assign high_exp__248 = 8'hff;
  assign is_result_nan__140 = eq_166708 & ne_166705 | eq_166710 & ne_166707 | has_pos_inf__68 & has_neg_inf__68;
  assign is_operand_inf__68 = eq_166708 & eq_166709 | eq_166710 & eq_166711;
  assign and_reduce_166943 = &wide_exponent__206[7:0];
  assign high_exp__320 = 8'hff;
  assign is_result_nan__12 = eq_166719 & ne_166716 | eq_166721 & ne_166718 | has_pos_inf__6 & has_neg_inf__6;
  assign is_operand_inf__6 = eq_166719 & eq_166720 | eq_166721 & eq_166722;
  assign and_reduce_166951 = &wide_exponent__18[7:0];
  assign fraction_shift__376 = 3'h3;
  assign fraction_shift__247 = 3'h4;
  assign is_subnormal__15 = $signed(exp__63) <= $signed(10'h000);
  assign high_exp__114 = 8'hff;
  assign result_exp__47 = is_result_nan__92 | has_inf_arg__47 | result_exp__46[8] | and_reduce_166841 ? high_exp__116 : result_exp__46[7:0];
  assign is_result_nan__63 = eq_166735 & ne_166732 | eq_166737 & ne_166734 | has_pos_inf__31 & has_neg_inf__31;
  assign is_operand_inf__31 = eq_166735 & eq_166736 | eq_166737 & eq_166738;
  assign and_reduce_166964 = &wide_exponent__93[7:0];
  assign fraction_shift__394 = 3'h3;
  assign fraction_shift__282 = 3'h4;
  assign is_subnormal__33 = $signed(exp__137) <= $signed(10'h000);
  assign high_exp__179 = 8'hff;
  assign result_exp__101 = is_result_nan__131 | has_inf_arg__67 | result_exp__99[8] | and_reduce_166853 ? high_exp__181 : result_exp__99[7:0];
  assign is_result_nan__102 = eq_166751 & ne_166748 | eq_166753 & ne_166750 | has_pos_inf__50 & has_neg_inf__50;
  assign is_operand_inf__50 = eq_166751 & eq_166752 | eq_166753 & eq_166754;
  assign and_reduce_166977 = &wide_exponent__150[7:0];
  assign fraction_shift__412 = 3'h3;
  assign fraction_shift__317 = 3'h4;
  assign is_subnormal__53 = $signed(exp__219) <= $signed(10'h000);
  assign high_exp__245 = 8'hff;
  assign result_exp__161 = is_result_nan__103 | has_inf_arg__53 | result_exp__159[8] | and_reduce_166867 ? high_exp__248 : result_exp__159[7:0];
  assign is_result_nan__141 = eq_166770 & ne_166767 | eq_166772 & ne_166769 | has_pos_inf__69 & has_neg_inf__69;
  assign is_operand_inf__69 = eq_166770 & eq_166771 | eq_166772 & eq_166773;
  assign and_reduce_166990 = &wide_exponent__207[7:0];
  assign fraction_shift__430 = 3'h3;
  assign fraction_shift__352 = 3'h4;
  assign is_subnormal__73 = $signed(exp__301) <= $signed(10'h000);
  assign high_exp__317 = 8'hff;
  assign result_exp__221 = is_result_nan__142 | has_inf_arg__73 | result_exp__219[8] | and_reduce_166881 ? high_exp__320 : result_exp__219[7:0];
  assign fraction_shift__377 = 3'h3;
  assign fraction_shift__248 = 3'h4;
  assign high_exp__115 = 8'hff;
  assign fraction_shift__45 = rounding_carry__14 ? fraction_shift__247 : fraction_shift__376;
  assign result_sign__439 = 1'h0;
  assign result_exponent__15 = is_result_nan__29 | is_operand_inf__14 | wide_exponent__44[8] | and_reduce_166895 ? high_exp__114 : wide_exponent__44[7:0];
  assign result_sign__440 = 1'h0;
  assign fraction_shift__395 = 3'h3;
  assign fraction_shift__283 = 3'h4;
  assign high_exp__180 = 8'hff;
  assign fraction_shift__92 = rounding_carry__30 ? fraction_shift__282 : fraction_shift__394;
  assign result_sign__536 = 1'h0;
  assign result_exponent__30 = is_result_nan__62 | is_operand_inf__30 | wide_exponent__92[8] | and_reduce_166911 ? high_exp__179 : wide_exponent__92[7:0];
  assign result_sign__537 = 1'h0;
  assign fraction_shift__413 = 3'h3;
  assign fraction_shift__318 = 3'h4;
  assign high_exp__246 = 8'hff;
  assign fraction_shift__149 = rounding_carry__49 ? fraction_shift__317 : fraction_shift__412;
  assign result_sign__636 = 1'h0;
  assign result_exponent__49 = is_result_nan__101 | is_operand_inf__49 | wide_exponent__149[8] | and_reduce_166927 ? high_exp__245 : wide_exponent__149[7:0];
  assign result_sign__637 = 1'h0;
  assign fraction_shift__431 = 3'h3;
  assign fraction_shift__353 = 3'h4;
  assign high_exp__318 = 8'hff;
  assign fraction_shift__206 = rounding_carry__68 ? fraction_shift__352 : fraction_shift__430;
  assign result_sign__744 = 1'h0;
  assign result_exponent__68 = is_result_nan__140 | is_operand_inf__68 | wide_exponent__206[8] | and_reduce_166943 ? high_exp__317 : wide_exponent__206[7:0];
  assign result_sign__745 = 1'h0;
  assign fraction_shift__18 = rounding_carry__6 ? fraction_shift__248 : fraction_shift__377;
  assign result_sign__441 = 1'h0;
  assign result_exponent__6 = is_result_nan__12 | is_operand_inf__6 | wide_exponent__18[8] | and_reduce_166951 ? high_exp__115 : wide_exponent__18[7:0];
  assign shrl_167050 = rounded_fraction__14 >> fraction_shift__45;
  assign concat_167054 = {result_sign__440, ~result_exp__47};
  assign fraction_shift__93 = rounding_carry__31 ? fraction_shift__283 : fraction_shift__395;
  assign result_sign__538 = 1'h0;
  assign result_exponent__31 = is_result_nan__63 | is_operand_inf__31 | wide_exponent__93[8] | and_reduce_166964 ? high_exp__180 : wide_exponent__93[7:0];
  assign shrl_167059 = rounded_fraction__30 >> fraction_shift__92;
  assign concat_167063 = {result_sign__537, ~result_exp__101};
  assign fraction_shift__150 = rounding_carry__50 ? fraction_shift__318 : fraction_shift__413;
  assign result_sign__638 = 1'h0;
  assign result_exponent__50 = is_result_nan__102 | is_operand_inf__50 | wide_exponent__150[8] | and_reduce_166977 ? high_exp__246 : wide_exponent__150[7:0];
  assign shrl_167068 = rounded_fraction__49 >> fraction_shift__149;
  assign concat_167072 = {result_sign__637, ~result_exp__161};
  assign fraction_shift__207 = rounding_carry__69 ? fraction_shift__353 : fraction_shift__431;
  assign result_sign__746 = 1'h0;
  assign result_exponent__69 = is_result_nan__141 | is_operand_inf__69 | wide_exponent__207[8] | and_reduce_166990 ? high_exp__318 : wide_exponent__207[7:0];
  assign shrl_167077 = rounded_fraction__68 >> fraction_shift__206;
  assign concat_167081 = {result_sign__745, ~result_exp__221};
  assign shrl_167082 = rounded_fraction__6 >> fraction_shift__18;
  assign result_fraction__87 = shrl_167050[22:0];
  assign result_fraction__90 = fraction__142[22:0];
  assign sum__15 = {result_sign__439, result_exponent__15} + concat_167054;
  assign shrl_167090 = rounded_fraction__31 >> fraction_shift__93;
  assign result_fraction__184 = shrl_167059[22:0];
  assign result_fraction__190 = fraction__302[22:0];
  assign sum__32 = {result_sign__536, result_exponent__30} + concat_167063;
  assign shrl_167098 = rounded_fraction__50 >> fraction_shift__150;
  assign result_fraction__301 = shrl_167068[22:0];
  assign result_fraction__307 = fraction__481[22:0];
  assign sum__51 = {result_sign__636, result_exponent__49} + concat_167072;
  assign shrl_167106 = rounded_fraction__69 >> fraction_shift__207;
  assign result_fraction__418 = shrl_167077[22:0];
  assign result_fraction__424 = fraction__660[22:0];
  assign sum__70 = {result_sign__744, result_exponent__68} + concat_167081;
  assign result_fraction__34 = shrl_167082[22:0];
  assign sum__7 = {result_sign__441, result_exponent__6} + concat_167054;
  assign result_fraction__88 = result_fraction__87 & {23{~(is_operand_inf__14 | wide_exponent__44[8] | and_reduce_166895 | ~((|wide_exponent__44[8:1]) | wide_exponent__44[0]))}};
  assign nan_fraction__93 = 23'h40_0000;
  assign result_fraction__91 = result_fraction__90 & {23{~(has_inf_arg__47 | result_exp__46[8] | and_reduce_166841 | is_subnormal__15)}};
  assign nan_fraction__95 = 23'h40_0000;
  assign result_fraction__185 = shrl_167090[22:0];
  assign sum__33 = {result_sign__538, result_exponent__31} + concat_167063;
  assign result_fraction__186 = result_fraction__184 & {23{~(is_operand_inf__30 | wide_exponent__92[8] | and_reduce_166911 | ~((|wide_exponent__92[8:1]) | wide_exponent__92[0]))}};
  assign nan_fraction__120 = 23'h40_0000;
  assign result_fraction__192 = result_fraction__190 & {23{~(has_inf_arg__67 | result_exp__99[8] | and_reduce_166853 | is_subnormal__33)}};
  assign nan_fraction__122 = 23'h40_0000;
  assign result_fraction__302 = shrl_167098[22:0];
  assign sum__52 = {result_sign__638, result_exponent__50} + concat_167072;
  assign result_fraction__303 = result_fraction__301 & {23{~(is_operand_inf__49 | wide_exponent__149[8] | and_reduce_166927 | ~((|wide_exponent__149[8:1]) | wide_exponent__149[0]))}};
  assign nan_fraction__148 = 23'h40_0000;
  assign result_fraction__309 = result_fraction__307 & {23{~(has_inf_arg__53 | result_exp__159[8] | and_reduce_166867 | is_subnormal__53)}};
  assign nan_fraction__150 = 23'h40_0000;
  assign result_fraction__419 = shrl_167106[22:0];
  assign sum__71 = {result_sign__746, result_exponent__69} + concat_167081;
  assign result_fraction__420 = result_fraction__418 & {23{~(is_operand_inf__68 | wide_exponent__206[8] | and_reduce_166943 | ~((|wide_exponent__206[8:1]) | wide_exponent__206[0]))}};
  assign nan_fraction__177 = 23'h40_0000;
  assign result_fraction__426 = result_fraction__424 & {23{~(has_inf_arg__73 | result_exp__219[8] | and_reduce_166881 | is_subnormal__73)}};
  assign nan_fraction__179 = 23'h40_0000;
  assign result_fraction__35 = result_fraction__34 & {23{~(is_operand_inf__6 | wide_exponent__18[8] | and_reduce_166951 | ~((|wide_exponent__18[8:1]) | wide_exponent__18[0]))}};
  assign nan_fraction__94 = 23'h40_0000;
  assign result_fraction__89 = is_result_nan__29 ? nan_fraction__93 : result_fraction__88;
  assign result_fraction__92 = is_result_nan__92 ? nan_fraction__95 : result_fraction__91;
  assign prod_bexp__62 = sum__15[8] ? result_exp__47 : result_exponent__15;
  assign x_bexp__762 = 8'h00;
  assign result_fraction__187 = result_fraction__185 & {23{~(is_operand_inf__31 | wide_exponent__93[8] | and_reduce_166964 | ~((|wide_exponent__93[8:1]) | wide_exponent__93[0]))}};
  assign nan_fraction__121 = 23'h40_0000;
  assign result_fraction__188 = is_result_nan__62 ? nan_fraction__120 : result_fraction__186;
  assign result_fraction__194 = is_result_nan__131 ? nan_fraction__122 : result_fraction__192;
  assign prod_bexp__123 = sum__32[8] ? result_exp__101 : result_exponent__30;
  assign x_bexp__763 = 8'h00;
  assign result_fraction__304 = result_fraction__302 & {23{~(is_operand_inf__50 | wide_exponent__150[8] | and_reduce_166977 | ~((|wide_exponent__150[8:1]) | wide_exponent__150[0]))}};
  assign nan_fraction__149 = 23'h40_0000;
  assign result_fraction__305 = is_result_nan__101 ? nan_fraction__148 : result_fraction__303;
  assign result_fraction__311 = is_result_nan__103 ? nan_fraction__150 : result_fraction__309;
  assign prod_bexp__195 = sum__51[8] ? result_exp__161 : result_exponent__49;
  assign x_bexp__764 = 8'h00;
  assign result_fraction__421 = result_fraction__419 & {23{~(is_operand_inf__69 | wide_exponent__207[8] | and_reduce_166990 | ~((|wide_exponent__207[8:1]) | wide_exponent__207[0]))}};
  assign nan_fraction__178 = 23'h40_0000;
  assign result_fraction__422 = is_result_nan__140 ? nan_fraction__177 : result_fraction__420;
  assign result_fraction__428 = is_result_nan__142 ? nan_fraction__179 : result_fraction__426;
  assign prod_bexp__267 = sum__70[8] ? result_exp__221 : result_exponent__68;
  assign x_bexp__765 = 8'h00;
  assign result_fraction__36 = is_result_nan__12 ? nan_fraction__94 : result_fraction__35;
  assign prod_bexp__26 = sum__7[8] ? result_exp__47 : result_exponent__6;
  assign x_bexp__766 = 8'h00;
  assign fraction_is_zero__14 = add_165914 == 26'h000_0000 & xddend_y__14[2:0] == 3'h0;
  assign prod_fraction__45 = sum__15[8] ? result_fraction__92 : result_fraction__89;
  assign incremented_sum__88 = sum__15[7:0] + 8'h01;
  assign result_fraction__189 = is_result_nan__63 ? nan_fraction__121 : result_fraction__187;
  assign prod_bexp__124 = sum__33[8] ? result_exp__101 : result_exponent__31;
  assign x_bexp__767 = 8'h00;
  assign fraction_is_zero__30 = add_165917 == 26'h000_0000 & xddend_y__29[2:0] == 3'h0;
  assign prod_fraction__91 = sum__32[8] ? result_fraction__194 : result_fraction__188;
  assign incremented_sum__106 = sum__32[7:0] + 8'h01;
  assign result_fraction__306 = is_result_nan__102 ? nan_fraction__149 : result_fraction__304;
  assign prod_bexp__196 = sum__52[8] ? result_exp__161 : result_exponent__50;
  assign x_bexp__768 = 8'h00;
  assign fraction_is_zero__49 = add_165920 == 26'h000_0000 & xddend_y__47[2:0] == 3'h0;
  assign prod_fraction__145 = sum__51[8] ? result_fraction__311 : result_fraction__305;
  assign incremented_sum__124 = sum__51[7:0] + 8'h01;
  assign result_fraction__423 = is_result_nan__141 ? nan_fraction__178 : result_fraction__421;
  assign prod_bexp__268 = sum__71[8] ? result_exp__221 : result_exponent__69;
  assign x_bexp__769 = 8'h00;
  assign fraction_is_zero__68 = add_165923 == 26'h000_0000 & xddend_y__65[2:0] == 3'h0;
  assign prod_fraction__199 = sum__70[8] ? result_fraction__428 : result_fraction__422;
  assign incremented_sum__142 = sum__70[7:0] + 8'h01;
  assign fraction_is_zero__6 = add_165924 == 26'h000_0000 & xddend_y__6[2:0] == 3'h0;
  assign prod_fraction__19 = sum__7[8] ? result_fraction__92 : result_fraction__36;
  assign incremented_sum__89 = sum__7[7:0] + 8'h01;
  assign wide_y__30 = {2'h1, prod_fraction__45, 3'h0};
  assign x_bexpbs_difference__16 = sum__15[8] ? incremented_sum__88 : ~sum__15[7:0];
  assign fraction_is_zero__31 = add_165927 == 26'h000_0000 & xddend_y__30[2:0] == 3'h0;
  assign prod_fraction__92 = sum__33[8] ? result_fraction__194 : result_fraction__189;
  assign incremented_sum__107 = sum__33[7:0] + 8'h01;
  assign wide_y__63 = {2'h1, prod_fraction__91, 3'h0};
  assign x_bexpbs_difference__31 = sum__32[8] ? incremented_sum__106 : ~sum__32[7:0];
  assign fraction_is_zero__50 = add_165930 == 26'h000_0000 & xddend_y__48[2:0] == 3'h0;
  assign prod_fraction__146 = sum__52[8] ? result_fraction__311 : result_fraction__306;
  assign incremented_sum__125 = sum__52[7:0] + 8'h01;
  assign wide_y__101 = {2'h1, prod_fraction__145, 3'h0};
  assign x_bexpbs_difference__49 = sum__51[8] ? incremented_sum__124 : ~sum__51[7:0];
  assign fraction_is_zero__69 = add_165933 == 26'h000_0000 & xddend_y__66[2:0] == 3'h0;
  assign prod_fraction__200 = sum__71[8] ? result_fraction__428 : result_fraction__423;
  assign incremented_sum__143 = sum__71[7:0] + 8'h01;
  assign wide_y__139 = {2'h1, prod_fraction__199, 3'h0};
  assign x_bexpbs_difference__67 = sum__70[8] ? incremented_sum__142 : ~sum__70[7:0];
  assign wide_y__13 = {2'h1, prod_fraction__19, 3'h0};
  assign x_bexpbs_difference__7 = sum__7[8] ? incremented_sum__89 : ~sum__7[7:0];
  assign concat_167315 = {~(add_165914[25] | fraction_is_zero__14), add_165914[25], fraction_is_zero__14};
  assign x_bexp__126 = sum__15[8] ? result_exponent__15 : result_exp__47;
  assign x_bexp__770 = 8'h00;
  assign wide_y__31 = wide_y__30 & {28{prod_bexp__62 != x_bexp__762}};
  assign sub_167321 = 8'h1c - x_bexpbs_difference__16;
  assign wide_y__64 = {2'h1, prod_fraction__92, 3'h0};
  assign x_bexpbs_difference__32 = sum__33[8] ? incremented_sum__107 : ~sum__33[7:0];
  assign concat_167327 = {~(add_165917[25] | fraction_is_zero__30), add_165917[25], fraction_is_zero__30};
  assign x_bexp__251 = sum__32[8] ? result_exponent__30 : result_exp__101;
  assign x_bexp__771 = 8'h00;
  assign wide_y__65 = wide_y__63 & {28{prod_bexp__123 != x_bexp__763}};
  assign sub_167333 = 8'h1c - x_bexpbs_difference__31;
  assign wide_y__102 = {2'h1, prod_fraction__146, 3'h0};
  assign x_bexpbs_difference__50 = sum__52[8] ? incremented_sum__125 : ~sum__52[7:0];
  assign concat_167339 = {~(add_165920[25] | fraction_is_zero__49), add_165920[25], fraction_is_zero__49};
  assign x_bexp__395 = sum__51[8] ? result_exponent__49 : result_exp__161;
  assign x_bexp__772 = 8'h00;
  assign wide_y__103 = wide_y__101 & {28{prod_bexp__195 != x_bexp__764}};
  assign sub_167345 = 8'h1c - x_bexpbs_difference__49;
  assign wide_y__140 = {2'h1, prod_fraction__200, 3'h0};
  assign x_bexpbs_difference__68 = sum__71[8] ? incremented_sum__143 : ~sum__71[7:0];
  assign concat_167351 = {~(add_165923[25] | fraction_is_zero__68), add_165923[25], fraction_is_zero__68};
  assign x_bexp__539 = sum__70[8] ? result_exponent__68 : result_exp__221;
  assign x_bexp__773 = 8'h00;
  assign wide_y__141 = wide_y__139 & {28{prod_bexp__267 != x_bexp__765}};
  assign sub_167357 = 8'h1c - x_bexpbs_difference__67;
  assign concat_167358 = {~(add_165924[25] | fraction_is_zero__6), add_165924[25], fraction_is_zero__6};
  assign x_bexp__54 = sum__7[8] ? result_exponent__6 : result_exp__47;
  assign x_bexp__774 = 8'h00;
  assign wide_y__14 = wide_y__13 & {28{prod_bexp__26 != x_bexp__766}};
  assign sub_167364 = 8'h1c - x_bexpbs_difference__7;
  assign result_sign__72 = x_sign__30 & prod_sign__14 & concat_167315[0] | ~prod_sign__14 & concat_167315[1] | prod_sign__14 & concat_167315[2];
  assign x_fraction__126 = sum__15[8] ? result_fraction__89 : result_fraction__92;
  assign dropped__15 = sub_167321 >= 8'h1c ? 28'h000_0000 : wide_y__31 << sub_167321;
  assign concat_167372 = {~(add_165927[25] | fraction_is_zero__31), add_165927[25], fraction_is_zero__31};
  assign x_bexp__252 = sum__33[8] ? result_exponent__31 : result_exp__101;
  assign x_bexp__775 = 8'h00;
  assign wide_y__66 = wide_y__64 & {28{prod_bexp__124 != x_bexp__767}};
  assign sub_167378 = 8'h1c - x_bexpbs_difference__32;
  assign result_sign__152 = x_sign__59 & prod_sign__29 & concat_167327[0] | ~prod_sign__29 & concat_167327[1] | prod_sign__29 & concat_167327[2];
  assign x_fraction__251 = sum__32[8] ? result_fraction__188 : result_fraction__194;
  assign dropped__32 = sub_167333 >= 8'h1c ? 28'h000_0000 : wide_y__65 << sub_167333;
  assign concat_167386 = {~(add_165930[25] | fraction_is_zero__50), add_165930[25], fraction_is_zero__50};
  assign x_bexp__396 = sum__52[8] ? result_exponent__50 : result_exp__161;
  assign x_bexp__776 = 8'h00;
  assign wide_y__104 = wide_y__102 & {28{prod_bexp__196 != x_bexp__768}};
  assign sub_167392 = 8'h1c - x_bexpbs_difference__50;
  assign result_sign__249 = x_sign__95 & prod_sign__47 & concat_167339[0] | ~prod_sign__47 & concat_167339[1] | prod_sign__47 & concat_167339[2];
  assign x_fraction__395 = sum__51[8] ? result_fraction__305 : result_fraction__311;
  assign dropped__51 = sub_167345 >= 8'h1c ? 28'h000_0000 : wide_y__103 << sub_167345;
  assign concat_167400 = {~(add_165933[25] | fraction_is_zero__69), add_165933[25], fraction_is_zero__69};
  assign x_bexp__540 = sum__71[8] ? result_exponent__69 : result_exp__221;
  assign x_bexp__777 = 8'h00;
  assign wide_y__142 = wide_y__140 & {28{prod_bexp__268 != x_bexp__769}};
  assign sub_167406 = 8'h1c - x_bexpbs_difference__68;
  assign result_sign__346 = x_sign__131 & prod_sign__65 & concat_167351[0] | ~prod_sign__65 & concat_167351[1] | prod_sign__65 & concat_167351[2];
  assign x_fraction__539 = sum__70[8] ? result_fraction__422 : result_fraction__428;
  assign dropped__70 = sub_167357 >= 8'h1c ? 28'h000_0000 : wide_y__141 << sub_167357;
  assign result_sign__28 = x_sign__12 & prod_sign__6 & concat_167358[0] | ~prod_sign__6 & concat_167358[1] | prod_sign__6 & concat_167358[2];
  assign x_fraction__54 = sum__7[8] ? result_fraction__36 : result_fraction__92;
  assign dropped__7 = sub_167364 >= 8'h1c ? 28'h000_0000 : wide_y__14 << sub_167364;
  assign result_sign__73 = is_operand_inf__14 ? ~has_pos_inf__14 : result_sign__72;
  assign wide_x__30 = {2'h1, x_fraction__126, 3'h0};
  assign result_sign__153 = x_sign__60 & prod_sign__30 & concat_167372[0] | ~prod_sign__30 & concat_167372[1] | prod_sign__30 & concat_167372[2];
  assign x_fraction__252 = sum__33[8] ? result_fraction__189 : result_fraction__194;
  assign dropped__33 = sub_167378 >= 8'h1c ? 28'h000_0000 : wide_y__66 << sub_167378;
  assign result_sign__154 = is_operand_inf__30 ? ~has_pos_inf__30 : result_sign__152;
  assign wide_x__63 = {2'h1, x_fraction__251, 3'h0};
  assign x_sign__98 = array_index_166097[31:31];
  assign result_sign__250 = x_sign__96 & prod_sign__48 & concat_167386[0] | ~prod_sign__48 & concat_167386[1] | prod_sign__48 & concat_167386[2];
  assign x_fraction__396 = sum__52[8] ? result_fraction__306 : result_fraction__311;
  assign dropped__52 = sub_167392 >= 8'h1c ? 28'h000_0000 : wide_y__104 << sub_167392;
  assign nand_167448 = ~(eq_166813 & ne_166814);
  assign result_sign__251 = is_operand_inf__49 ? ~has_pos_inf__49 : result_sign__249;
  assign wide_x__101 = {2'h1, x_fraction__395, 3'h0};
  assign x_sign__134 = array_index_166111[31:31];
  assign result_sign__347 = x_sign__132 & prod_sign__66 & concat_167400[0] | ~prod_sign__66 & concat_167400[1] | prod_sign__66 & concat_167400[2];
  assign x_fraction__540 = sum__71[8] ? result_fraction__423 : result_fraction__428;
  assign dropped__71 = sub_167406 >= 8'h1c ? 28'h000_0000 : wide_y__142 << sub_167406;
  assign nand_167463 = ~(is_result_nan__108 & ne_166827);
  assign result_sign__348 = is_operand_inf__68 ? ~has_pos_inf__68 : result_sign__346;
  assign wide_x__139 = {2'h1, x_fraction__539, 3'h0};
  assign result_sign__29 = is_operand_inf__6 ? ~has_pos_inf__6 : result_sign__28;
  assign wide_x__13 = {2'h1, x_fraction__54, 3'h0};
  assign result_sign__76 = nand_162587 & x_sign__86;
  assign result_sign__74 = ~is_result_nan__29 & result_sign__73;
  assign wide_x__31 = wide_x__30 & {28{x_bexp__126 != x_bexp__770}};
  assign result_sign__155 = is_operand_inf__31 ? ~has_pos_inf__31 : result_sign__153;
  assign wide_x__64 = {2'h1, x_fraction__252, 3'h0};
  assign result_sign__160 = nand_162600 & x_sign__122;
  assign result_sign__156 = ~is_result_nan__62 & result_sign__154;
  assign wide_x__65 = wide_x__63 & {28{x_bexp__251 != x_bexp__771}};
  assign result_sign__256 = ~x_sign__98;
  assign result_sign__252 = is_operand_inf__50 ? ~has_pos_inf__50 : result_sign__250;
  assign wide_x__102 = {2'h1, x_fraction__396, 3'h0};
  assign result_sign__257 = nand_167448 & x_sign__98;
  assign result_sign__253 = ~is_result_nan__101 & result_sign__251;
  assign wide_x__103 = wide_x__101 & {28{x_bexp__395 != x_bexp__772}};
  assign result_sign__353 = ~x_sign__134;
  assign result_sign__349 = is_operand_inf__69 ? ~has_pos_inf__69 : result_sign__347;
  assign wide_x__140 = {2'h1, x_fraction__540, 3'h0};
  assign result_sign__354 = nand_167463 & x_sign__134;
  assign result_sign__350 = ~is_result_nan__140 & result_sign__348;
  assign wide_x__141 = wide_x__139 & {28{x_bexp__539 != x_bexp__773}};
  assign result_sign__30 = ~is_result_nan__12 & result_sign__29;
  assign wide_x__14 = wide_x__13 & {28{x_bexp__54 != x_bexp__774}};
  assign x_sign__32 = sum__15[8] ? result_sign__74 : result_sign__76;
  assign prod_sign__15 = sum__15[8] ? result_sign__76 : result_sign__74;
  assign neg_167522 = -wide_x__31;
  assign sticky__47 = {27'h000_0000, dropped__15[27:3] != 25'h000_0000};
  assign result_sign__157 = ~is_result_nan__63 & result_sign__155;
  assign wide_x__66 = wide_x__64 & {28{x_bexp__252 != x_bexp__775}};
  assign x_sign__63 = sum__32[8] ? result_sign__156 : result_sign__160;
  assign prod_sign__31 = sum__32[8] ? result_sign__160 : result_sign__156;
  assign neg_167531 = -wide_x__65;
  assign sticky__100 = {27'h000_0000, dropped__32[27:3] != 25'h000_0000};
  assign result_sign__258 = nand_167448 & result_sign__256;
  assign result_sign__254 = ~is_result_nan__102 & result_sign__252;
  assign wide_x__104 = wide_x__102 & {28{x_bexp__396 != x_bexp__776}};
  assign x_sign__99 = sum__51[8] ? result_sign__253 : result_sign__257;
  assign prod_sign__49 = sum__51[8] ? result_sign__257 : result_sign__253;
  assign neg_167541 = -wide_x__103;
  assign sticky__159 = {27'h000_0000, dropped__51[27:3] != 25'h000_0000};
  assign result_sign__355 = nand_167463 & result_sign__353;
  assign result_sign__351 = ~is_result_nan__141 & result_sign__349;
  assign wide_x__142 = wide_x__140 & {28{x_bexp__540 != x_bexp__777}};
  assign x_sign__135 = sum__70[8] ? result_sign__350 : result_sign__354;
  assign prod_sign__67 = sum__70[8] ? result_sign__354 : result_sign__350;
  assign neg_167551 = -wide_x__141;
  assign sticky__218 = {27'h000_0000, dropped__70[27:3] != 25'h000_0000};
  assign x_sign__14 = sum__7[8] ? result_sign__30 : result_sign__228;
  assign prod_sign__7 = sum__7[8] ? result_sign__228 : result_sign__30;
  assign neg_167556 = -wide_x__14;
  assign sticky__21 = {27'h000_0000, dropped__7[27:3] != 25'h000_0000};
  assign xddend_y__15 = (x_bexpbs_difference__16 >= 8'h1c ? 28'h000_0000 : wide_y__31 >> x_bexpbs_difference__16) | sticky__47;
  assign x_sign__64 = sum__33[8] ? result_sign__157 : result_sign__325;
  assign prod_sign__32 = sum__33[8] ? result_sign__325 : result_sign__157;
  assign neg_167565 = -wide_x__66;
  assign sticky__101 = {27'h000_0000, dropped__33[27:3] != 25'h000_0000};
  assign xddend_y__31 = (x_bexpbs_difference__31 >= 8'h1c ? 28'h000_0000 : wide_y__65 >> x_bexpbs_difference__31) | sticky__100;
  assign x_sign__100 = sum__52[8] ? result_sign__254 : result_sign__258;
  assign prod_sign__50 = sum__52[8] ? result_sign__258 : result_sign__254;
  assign neg_167574 = -wide_x__104;
  assign sticky__160 = {27'h000_0000, dropped__52[27:3] != 25'h000_0000};
  assign xddend_y__49 = (x_bexpbs_difference__49 >= 8'h1c ? 28'h000_0000 : wide_y__103 >> x_bexpbs_difference__49) | sticky__159;
  assign x_sign__136 = sum__71[8] ? result_sign__351 : result_sign__355;
  assign prod_sign__68 = sum__71[8] ? result_sign__355 : result_sign__351;
  assign neg_167583 = -wide_x__142;
  assign sticky__219 = {27'h000_0000, dropped__71[27:3] != 25'h000_0000};
  assign xddend_y__67 = (x_bexpbs_difference__67 >= 8'h1c ? 28'h000_0000 : wide_y__141 >> x_bexpbs_difference__67) | sticky__218;
  assign xddend_y__7 = (x_bexpbs_difference__7 >= 8'h1c ? 28'h000_0000 : wide_y__14 >> x_bexpbs_difference__7) | sticky__21;
  assign sel_167594 = x_sign__32 ^ prod_sign__15 ? neg_167522[27:3] : wide_x__31[27:3];
  assign result_sign__1050 = 1'h0;
  assign xddend_y__32 = (x_bexpbs_difference__32 >= 8'h1c ? 28'h000_0000 : wide_y__66 >> x_bexpbs_difference__32) | sticky__101;
  assign sel_167601 = x_sign__63 ^ prod_sign__31 ? neg_167531[27:3] : wide_x__65[27:3];
  assign result_sign__1051 = 1'h0;
  assign xddend_y__50 = (x_bexpbs_difference__50 >= 8'h1c ? 28'h000_0000 : wide_y__104 >> x_bexpbs_difference__50) | sticky__160;
  assign sel_167608 = x_sign__99 ^ prod_sign__49 ? neg_167541[27:3] : wide_x__103[27:3];
  assign result_sign__1052 = 1'h0;
  assign xddend_y__68 = (x_bexpbs_difference__68 >= 8'h1c ? 28'h000_0000 : wide_y__142 >> x_bexpbs_difference__68) | sticky__219;
  assign sel_167615 = x_sign__135 ^ prod_sign__67 ? neg_167551[27:3] : wide_x__141[27:3];
  assign result_sign__1053 = 1'h0;
  assign sel_167618 = x_sign__14 ^ prod_sign__7 ? neg_167556[27:3] : wide_x__14[27:3];
  assign result_sign__1054 = 1'h0;
  assign sel_167623 = x_sign__64 ^ prod_sign__32 ? neg_167565[27:3] : wide_x__66[27:3];
  assign result_sign__1055 = 1'h0;
  assign sel_167628 = x_sign__100 ^ prod_sign__50 ? neg_167574[27:3] : wide_x__104[27:3];
  assign result_sign__1056 = 1'h0;
  assign sel_167633 = x_sign__136 ^ prod_sign__68 ? neg_167583[27:3] : wide_x__142[27:3];
  assign result_sign__1057 = 1'h0;
  assign add_167640 = {{1{sel_167594[24]}}, sel_167594} + {result_sign__1050, xddend_y__15[27:3]};
  assign add_167643 = {{1{sel_167601[24]}}, sel_167601} + {result_sign__1051, xddend_y__31[27:3]};
  assign add_167646 = {{1{sel_167608[24]}}, sel_167608} + {result_sign__1052, xddend_y__49[27:3]};
  assign add_167649 = {{1{sel_167615[24]}}, sel_167615} + {result_sign__1053, xddend_y__67[27:3]};
  assign add_167650 = {{1{sel_167618[24]}}, sel_167618} + {result_sign__1054, xddend_y__7[27:3]};
  assign add_167653 = {{1{sel_167623[24]}}, sel_167623} + {result_sign__1055, xddend_y__32[27:3]};
  assign add_167656 = {{1{sel_167628[24]}}, sel_167628} + {result_sign__1056, xddend_y__50[27:3]};
  assign add_167659 = {{1{sel_167633[24]}}, sel_167633} + {result_sign__1057, xddend_y__68[27:3]};
  assign concat_167664 = {add_167640[24:0], xddend_y__15[2:0]};
  assign concat_167667 = {add_167643[24:0], xddend_y__31[2:0]};
  assign concat_167670 = {add_167646[24:0], xddend_y__49[2:0]};
  assign concat_167673 = {add_167649[24:0], xddend_y__67[2:0]};
  assign concat_167674 = {add_167650[24:0], xddend_y__7[2:0]};
  assign concat_167677 = {add_167653[24:0], xddend_y__32[2:0]};
  assign concat_167680 = {add_167656[24:0], xddend_y__50[2:0]};
  assign concat_167683 = {add_167659[24:0], xddend_y__68[2:0]};
  assign xbs_fraction__15 = add_167640[25] ? -concat_167664 : concat_167664;
  assign xbs_fraction__31 = add_167643[25] ? -concat_167667 : concat_167667;
  assign xbs_fraction__49 = add_167646[25] ? -concat_167670 : concat_167670;
  assign xbs_fraction__67 = add_167649[25] ? -concat_167673 : concat_167673;
  assign xbs_fraction__7 = add_167650[25] ? -concat_167674 : concat_167674;
  assign reverse_167699 = {xbs_fraction__15[0], xbs_fraction__15[1], xbs_fraction__15[2], xbs_fraction__15[3], xbs_fraction__15[4], xbs_fraction__15[5], xbs_fraction__15[6], xbs_fraction__15[7], xbs_fraction__15[8], xbs_fraction__15[9], xbs_fraction__15[10], xbs_fraction__15[11], xbs_fraction__15[12], xbs_fraction__15[13], xbs_fraction__15[14], xbs_fraction__15[15], xbs_fraction__15[16], xbs_fraction__15[17], xbs_fraction__15[18], xbs_fraction__15[19], xbs_fraction__15[20], xbs_fraction__15[21], xbs_fraction__15[22], xbs_fraction__15[23], xbs_fraction__15[24], xbs_fraction__15[25], xbs_fraction__15[26], xbs_fraction__15[27]};
  assign xbs_fraction__32 = add_167653[25] ? -concat_167677 : concat_167677;
  assign reverse_167701 = {xbs_fraction__31[0], xbs_fraction__31[1], xbs_fraction__31[2], xbs_fraction__31[3], xbs_fraction__31[4], xbs_fraction__31[5], xbs_fraction__31[6], xbs_fraction__31[7], xbs_fraction__31[8], xbs_fraction__31[9], xbs_fraction__31[10], xbs_fraction__31[11], xbs_fraction__31[12], xbs_fraction__31[13], xbs_fraction__31[14], xbs_fraction__31[15], xbs_fraction__31[16], xbs_fraction__31[17], xbs_fraction__31[18], xbs_fraction__31[19], xbs_fraction__31[20], xbs_fraction__31[21], xbs_fraction__31[22], xbs_fraction__31[23], xbs_fraction__31[24], xbs_fraction__31[25], xbs_fraction__31[26], xbs_fraction__31[27]};
  assign xbs_fraction__50 = add_167656[25] ? -concat_167680 : concat_167680;
  assign reverse_167703 = {xbs_fraction__49[0], xbs_fraction__49[1], xbs_fraction__49[2], xbs_fraction__49[3], xbs_fraction__49[4], xbs_fraction__49[5], xbs_fraction__49[6], xbs_fraction__49[7], xbs_fraction__49[8], xbs_fraction__49[9], xbs_fraction__49[10], xbs_fraction__49[11], xbs_fraction__49[12], xbs_fraction__49[13], xbs_fraction__49[14], xbs_fraction__49[15], xbs_fraction__49[16], xbs_fraction__49[17], xbs_fraction__49[18], xbs_fraction__49[19], xbs_fraction__49[20], xbs_fraction__49[21], xbs_fraction__49[22], xbs_fraction__49[23], xbs_fraction__49[24], xbs_fraction__49[25], xbs_fraction__49[26], xbs_fraction__49[27]};
  assign xbs_fraction__68 = add_167659[25] ? -concat_167683 : concat_167683;
  assign reverse_167705 = {xbs_fraction__67[0], xbs_fraction__67[1], xbs_fraction__67[2], xbs_fraction__67[3], xbs_fraction__67[4], xbs_fraction__67[5], xbs_fraction__67[6], xbs_fraction__67[7], xbs_fraction__67[8], xbs_fraction__67[9], xbs_fraction__67[10], xbs_fraction__67[11], xbs_fraction__67[12], xbs_fraction__67[13], xbs_fraction__67[14], xbs_fraction__67[15], xbs_fraction__67[16], xbs_fraction__67[17], xbs_fraction__67[18], xbs_fraction__67[19], xbs_fraction__67[20], xbs_fraction__67[21], xbs_fraction__67[22], xbs_fraction__67[23], xbs_fraction__67[24], xbs_fraction__67[25], xbs_fraction__67[26], xbs_fraction__67[27]};
  assign reverse_167706 = {xbs_fraction__7[0], xbs_fraction__7[1], xbs_fraction__7[2], xbs_fraction__7[3], xbs_fraction__7[4], xbs_fraction__7[5], xbs_fraction__7[6], xbs_fraction__7[7], xbs_fraction__7[8], xbs_fraction__7[9], xbs_fraction__7[10], xbs_fraction__7[11], xbs_fraction__7[12], xbs_fraction__7[13], xbs_fraction__7[14], xbs_fraction__7[15], xbs_fraction__7[16], xbs_fraction__7[17], xbs_fraction__7[18], xbs_fraction__7[19], xbs_fraction__7[20], xbs_fraction__7[21], xbs_fraction__7[22], xbs_fraction__7[23], xbs_fraction__7[24], xbs_fraction__7[25], xbs_fraction__7[26], xbs_fraction__7[27]};
  assign one_hot_167707 = {reverse_167699[27:0] == 28'h000_0000, reverse_167699[27] && reverse_167699[26:0] == 27'h000_0000, reverse_167699[26] && reverse_167699[25:0] == 26'h000_0000, reverse_167699[25] && reverse_167699[24:0] == 25'h000_0000, reverse_167699[24] && reverse_167699[23:0] == 24'h00_0000, reverse_167699[23] && reverse_167699[22:0] == 23'h00_0000, reverse_167699[22] && reverse_167699[21:0] == 22'h00_0000, reverse_167699[21] && reverse_167699[20:0] == 21'h00_0000, reverse_167699[20] && reverse_167699[19:0] == 20'h0_0000, reverse_167699[19] && reverse_167699[18:0] == 19'h0_0000, reverse_167699[18] && reverse_167699[17:0] == 18'h0_0000, reverse_167699[17] && reverse_167699[16:0] == 17'h0_0000, reverse_167699[16] && reverse_167699[15:0] == 16'h0000, reverse_167699[15] && reverse_167699[14:0] == 15'h0000, reverse_167699[14] && reverse_167699[13:0] == 14'h0000, reverse_167699[13] && reverse_167699[12:0] == 13'h0000, reverse_167699[12] && reverse_167699[11:0] == 12'h000, reverse_167699[11] && reverse_167699[10:0] == 11'h000, reverse_167699[10] && reverse_167699[9:0] == 10'h000, reverse_167699[9] && reverse_167699[8:0] == 9'h000, reverse_167699[8] && reverse_167699[7:0] == 8'h00, reverse_167699[7] && reverse_167699[6:0] == 7'h00, reverse_167699[6] && reverse_167699[5:0] == 6'h00, reverse_167699[5] && reverse_167699[4:0] == 5'h00, reverse_167699[4] && reverse_167699[3:0] == 4'h0, reverse_167699[3] && reverse_167699[2:0] == 3'h0, reverse_167699[2] && reverse_167699[1:0] == 2'h0, reverse_167699[1] && !reverse_167699[0], reverse_167699[0]};
  assign reverse_167708 = {xbs_fraction__32[0], xbs_fraction__32[1], xbs_fraction__32[2], xbs_fraction__32[3], xbs_fraction__32[4], xbs_fraction__32[5], xbs_fraction__32[6], xbs_fraction__32[7], xbs_fraction__32[8], xbs_fraction__32[9], xbs_fraction__32[10], xbs_fraction__32[11], xbs_fraction__32[12], xbs_fraction__32[13], xbs_fraction__32[14], xbs_fraction__32[15], xbs_fraction__32[16], xbs_fraction__32[17], xbs_fraction__32[18], xbs_fraction__32[19], xbs_fraction__32[20], xbs_fraction__32[21], xbs_fraction__32[22], xbs_fraction__32[23], xbs_fraction__32[24], xbs_fraction__32[25], xbs_fraction__32[26], xbs_fraction__32[27]};
  assign one_hot_167709 = {reverse_167701[27:0] == 28'h000_0000, reverse_167701[27] && reverse_167701[26:0] == 27'h000_0000, reverse_167701[26] && reverse_167701[25:0] == 26'h000_0000, reverse_167701[25] && reverse_167701[24:0] == 25'h000_0000, reverse_167701[24] && reverse_167701[23:0] == 24'h00_0000, reverse_167701[23] && reverse_167701[22:0] == 23'h00_0000, reverse_167701[22] && reverse_167701[21:0] == 22'h00_0000, reverse_167701[21] && reverse_167701[20:0] == 21'h00_0000, reverse_167701[20] && reverse_167701[19:0] == 20'h0_0000, reverse_167701[19] && reverse_167701[18:0] == 19'h0_0000, reverse_167701[18] && reverse_167701[17:0] == 18'h0_0000, reverse_167701[17] && reverse_167701[16:0] == 17'h0_0000, reverse_167701[16] && reverse_167701[15:0] == 16'h0000, reverse_167701[15] && reverse_167701[14:0] == 15'h0000, reverse_167701[14] && reverse_167701[13:0] == 14'h0000, reverse_167701[13] && reverse_167701[12:0] == 13'h0000, reverse_167701[12] && reverse_167701[11:0] == 12'h000, reverse_167701[11] && reverse_167701[10:0] == 11'h000, reverse_167701[10] && reverse_167701[9:0] == 10'h000, reverse_167701[9] && reverse_167701[8:0] == 9'h000, reverse_167701[8] && reverse_167701[7:0] == 8'h00, reverse_167701[7] && reverse_167701[6:0] == 7'h00, reverse_167701[6] && reverse_167701[5:0] == 6'h00, reverse_167701[5] && reverse_167701[4:0] == 5'h00, reverse_167701[4] && reverse_167701[3:0] == 4'h0, reverse_167701[3] && reverse_167701[2:0] == 3'h0, reverse_167701[2] && reverse_167701[1:0] == 2'h0, reverse_167701[1] && !reverse_167701[0], reverse_167701[0]};
  assign reverse_167710 = {xbs_fraction__50[0], xbs_fraction__50[1], xbs_fraction__50[2], xbs_fraction__50[3], xbs_fraction__50[4], xbs_fraction__50[5], xbs_fraction__50[6], xbs_fraction__50[7], xbs_fraction__50[8], xbs_fraction__50[9], xbs_fraction__50[10], xbs_fraction__50[11], xbs_fraction__50[12], xbs_fraction__50[13], xbs_fraction__50[14], xbs_fraction__50[15], xbs_fraction__50[16], xbs_fraction__50[17], xbs_fraction__50[18], xbs_fraction__50[19], xbs_fraction__50[20], xbs_fraction__50[21], xbs_fraction__50[22], xbs_fraction__50[23], xbs_fraction__50[24], xbs_fraction__50[25], xbs_fraction__50[26], xbs_fraction__50[27]};
  assign one_hot_167711 = {reverse_167703[27:0] == 28'h000_0000, reverse_167703[27] && reverse_167703[26:0] == 27'h000_0000, reverse_167703[26] && reverse_167703[25:0] == 26'h000_0000, reverse_167703[25] && reverse_167703[24:0] == 25'h000_0000, reverse_167703[24] && reverse_167703[23:0] == 24'h00_0000, reverse_167703[23] && reverse_167703[22:0] == 23'h00_0000, reverse_167703[22] && reverse_167703[21:0] == 22'h00_0000, reverse_167703[21] && reverse_167703[20:0] == 21'h00_0000, reverse_167703[20] && reverse_167703[19:0] == 20'h0_0000, reverse_167703[19] && reverse_167703[18:0] == 19'h0_0000, reverse_167703[18] && reverse_167703[17:0] == 18'h0_0000, reverse_167703[17] && reverse_167703[16:0] == 17'h0_0000, reverse_167703[16] && reverse_167703[15:0] == 16'h0000, reverse_167703[15] && reverse_167703[14:0] == 15'h0000, reverse_167703[14] && reverse_167703[13:0] == 14'h0000, reverse_167703[13] && reverse_167703[12:0] == 13'h0000, reverse_167703[12] && reverse_167703[11:0] == 12'h000, reverse_167703[11] && reverse_167703[10:0] == 11'h000, reverse_167703[10] && reverse_167703[9:0] == 10'h000, reverse_167703[9] && reverse_167703[8:0] == 9'h000, reverse_167703[8] && reverse_167703[7:0] == 8'h00, reverse_167703[7] && reverse_167703[6:0] == 7'h00, reverse_167703[6] && reverse_167703[5:0] == 6'h00, reverse_167703[5] && reverse_167703[4:0] == 5'h00, reverse_167703[4] && reverse_167703[3:0] == 4'h0, reverse_167703[3] && reverse_167703[2:0] == 3'h0, reverse_167703[2] && reverse_167703[1:0] == 2'h0, reverse_167703[1] && !reverse_167703[0], reverse_167703[0]};
  assign reverse_167712 = {xbs_fraction__68[0], xbs_fraction__68[1], xbs_fraction__68[2], xbs_fraction__68[3], xbs_fraction__68[4], xbs_fraction__68[5], xbs_fraction__68[6], xbs_fraction__68[7], xbs_fraction__68[8], xbs_fraction__68[9], xbs_fraction__68[10], xbs_fraction__68[11], xbs_fraction__68[12], xbs_fraction__68[13], xbs_fraction__68[14], xbs_fraction__68[15], xbs_fraction__68[16], xbs_fraction__68[17], xbs_fraction__68[18], xbs_fraction__68[19], xbs_fraction__68[20], xbs_fraction__68[21], xbs_fraction__68[22], xbs_fraction__68[23], xbs_fraction__68[24], xbs_fraction__68[25], xbs_fraction__68[26], xbs_fraction__68[27]};
  assign one_hot_167713 = {reverse_167705[27:0] == 28'h000_0000, reverse_167705[27] && reverse_167705[26:0] == 27'h000_0000, reverse_167705[26] && reverse_167705[25:0] == 26'h000_0000, reverse_167705[25] && reverse_167705[24:0] == 25'h000_0000, reverse_167705[24] && reverse_167705[23:0] == 24'h00_0000, reverse_167705[23] && reverse_167705[22:0] == 23'h00_0000, reverse_167705[22] && reverse_167705[21:0] == 22'h00_0000, reverse_167705[21] && reverse_167705[20:0] == 21'h00_0000, reverse_167705[20] && reverse_167705[19:0] == 20'h0_0000, reverse_167705[19] && reverse_167705[18:0] == 19'h0_0000, reverse_167705[18] && reverse_167705[17:0] == 18'h0_0000, reverse_167705[17] && reverse_167705[16:0] == 17'h0_0000, reverse_167705[16] && reverse_167705[15:0] == 16'h0000, reverse_167705[15] && reverse_167705[14:0] == 15'h0000, reverse_167705[14] && reverse_167705[13:0] == 14'h0000, reverse_167705[13] && reverse_167705[12:0] == 13'h0000, reverse_167705[12] && reverse_167705[11:0] == 12'h000, reverse_167705[11] && reverse_167705[10:0] == 11'h000, reverse_167705[10] && reverse_167705[9:0] == 10'h000, reverse_167705[9] && reverse_167705[8:0] == 9'h000, reverse_167705[8] && reverse_167705[7:0] == 8'h00, reverse_167705[7] && reverse_167705[6:0] == 7'h00, reverse_167705[6] && reverse_167705[5:0] == 6'h00, reverse_167705[5] && reverse_167705[4:0] == 5'h00, reverse_167705[4] && reverse_167705[3:0] == 4'h0, reverse_167705[3] && reverse_167705[2:0] == 3'h0, reverse_167705[2] && reverse_167705[1:0] == 2'h0, reverse_167705[1] && !reverse_167705[0], reverse_167705[0]};
  assign one_hot_167714 = {reverse_167706[27:0] == 28'h000_0000, reverse_167706[27] && reverse_167706[26:0] == 27'h000_0000, reverse_167706[26] && reverse_167706[25:0] == 26'h000_0000, reverse_167706[25] && reverse_167706[24:0] == 25'h000_0000, reverse_167706[24] && reverse_167706[23:0] == 24'h00_0000, reverse_167706[23] && reverse_167706[22:0] == 23'h00_0000, reverse_167706[22] && reverse_167706[21:0] == 22'h00_0000, reverse_167706[21] && reverse_167706[20:0] == 21'h00_0000, reverse_167706[20] && reverse_167706[19:0] == 20'h0_0000, reverse_167706[19] && reverse_167706[18:0] == 19'h0_0000, reverse_167706[18] && reverse_167706[17:0] == 18'h0_0000, reverse_167706[17] && reverse_167706[16:0] == 17'h0_0000, reverse_167706[16] && reverse_167706[15:0] == 16'h0000, reverse_167706[15] && reverse_167706[14:0] == 15'h0000, reverse_167706[14] && reverse_167706[13:0] == 14'h0000, reverse_167706[13] && reverse_167706[12:0] == 13'h0000, reverse_167706[12] && reverse_167706[11:0] == 12'h000, reverse_167706[11] && reverse_167706[10:0] == 11'h000, reverse_167706[10] && reverse_167706[9:0] == 10'h000, reverse_167706[9] && reverse_167706[8:0] == 9'h000, reverse_167706[8] && reverse_167706[7:0] == 8'h00, reverse_167706[7] && reverse_167706[6:0] == 7'h00, reverse_167706[6] && reverse_167706[5:0] == 6'h00, reverse_167706[5] && reverse_167706[4:0] == 5'h00, reverse_167706[4] && reverse_167706[3:0] == 4'h0, reverse_167706[3] && reverse_167706[2:0] == 3'h0, reverse_167706[2] && reverse_167706[1:0] == 2'h0, reverse_167706[1] && !reverse_167706[0], reverse_167706[0]};
  assign encode_167715 = {one_hot_167707[16] | one_hot_167707[17] | one_hot_167707[18] | one_hot_167707[19] | one_hot_167707[20] | one_hot_167707[21] | one_hot_167707[22] | one_hot_167707[23] | one_hot_167707[24] | one_hot_167707[25] | one_hot_167707[26] | one_hot_167707[27] | one_hot_167707[28], one_hot_167707[8] | one_hot_167707[9] | one_hot_167707[10] | one_hot_167707[11] | one_hot_167707[12] | one_hot_167707[13] | one_hot_167707[14] | one_hot_167707[15] | one_hot_167707[24] | one_hot_167707[25] | one_hot_167707[26] | one_hot_167707[27] | one_hot_167707[28], one_hot_167707[4] | one_hot_167707[5] | one_hot_167707[6] | one_hot_167707[7] | one_hot_167707[12] | one_hot_167707[13] | one_hot_167707[14] | one_hot_167707[15] | one_hot_167707[20] | one_hot_167707[21] | one_hot_167707[22] | one_hot_167707[23] | one_hot_167707[28], one_hot_167707[2] | one_hot_167707[3] | one_hot_167707[6] | one_hot_167707[7] | one_hot_167707[10] | one_hot_167707[11] | one_hot_167707[14] | one_hot_167707[15] | one_hot_167707[18] | one_hot_167707[19] | one_hot_167707[22] | one_hot_167707[23] | one_hot_167707[26] | one_hot_167707[27], one_hot_167707[1] | one_hot_167707[3] | one_hot_167707[5] | one_hot_167707[7] | one_hot_167707[9] | one_hot_167707[11] | one_hot_167707[13] | one_hot_167707[15] | one_hot_167707[17] | one_hot_167707[19] | one_hot_167707[21] | one_hot_167707[23] | one_hot_167707[25] | one_hot_167707[27]};
  assign one_hot_167716 = {reverse_167708[27:0] == 28'h000_0000, reverse_167708[27] && reverse_167708[26:0] == 27'h000_0000, reverse_167708[26] && reverse_167708[25:0] == 26'h000_0000, reverse_167708[25] && reverse_167708[24:0] == 25'h000_0000, reverse_167708[24] && reverse_167708[23:0] == 24'h00_0000, reverse_167708[23] && reverse_167708[22:0] == 23'h00_0000, reverse_167708[22] && reverse_167708[21:0] == 22'h00_0000, reverse_167708[21] && reverse_167708[20:0] == 21'h00_0000, reverse_167708[20] && reverse_167708[19:0] == 20'h0_0000, reverse_167708[19] && reverse_167708[18:0] == 19'h0_0000, reverse_167708[18] && reverse_167708[17:0] == 18'h0_0000, reverse_167708[17] && reverse_167708[16:0] == 17'h0_0000, reverse_167708[16] && reverse_167708[15:0] == 16'h0000, reverse_167708[15] && reverse_167708[14:0] == 15'h0000, reverse_167708[14] && reverse_167708[13:0] == 14'h0000, reverse_167708[13] && reverse_167708[12:0] == 13'h0000, reverse_167708[12] && reverse_167708[11:0] == 12'h000, reverse_167708[11] && reverse_167708[10:0] == 11'h000, reverse_167708[10] && reverse_167708[9:0] == 10'h000, reverse_167708[9] && reverse_167708[8:0] == 9'h000, reverse_167708[8] && reverse_167708[7:0] == 8'h00, reverse_167708[7] && reverse_167708[6:0] == 7'h00, reverse_167708[6] && reverse_167708[5:0] == 6'h00, reverse_167708[5] && reverse_167708[4:0] == 5'h00, reverse_167708[4] && reverse_167708[3:0] == 4'h0, reverse_167708[3] && reverse_167708[2:0] == 3'h0, reverse_167708[2] && reverse_167708[1:0] == 2'h0, reverse_167708[1] && !reverse_167708[0], reverse_167708[0]};
  assign encode_167717 = {one_hot_167709[16] | one_hot_167709[17] | one_hot_167709[18] | one_hot_167709[19] | one_hot_167709[20] | one_hot_167709[21] | one_hot_167709[22] | one_hot_167709[23] | one_hot_167709[24] | one_hot_167709[25] | one_hot_167709[26] | one_hot_167709[27] | one_hot_167709[28], one_hot_167709[8] | one_hot_167709[9] | one_hot_167709[10] | one_hot_167709[11] | one_hot_167709[12] | one_hot_167709[13] | one_hot_167709[14] | one_hot_167709[15] | one_hot_167709[24] | one_hot_167709[25] | one_hot_167709[26] | one_hot_167709[27] | one_hot_167709[28], one_hot_167709[4] | one_hot_167709[5] | one_hot_167709[6] | one_hot_167709[7] | one_hot_167709[12] | one_hot_167709[13] | one_hot_167709[14] | one_hot_167709[15] | one_hot_167709[20] | one_hot_167709[21] | one_hot_167709[22] | one_hot_167709[23] | one_hot_167709[28], one_hot_167709[2] | one_hot_167709[3] | one_hot_167709[6] | one_hot_167709[7] | one_hot_167709[10] | one_hot_167709[11] | one_hot_167709[14] | one_hot_167709[15] | one_hot_167709[18] | one_hot_167709[19] | one_hot_167709[22] | one_hot_167709[23] | one_hot_167709[26] | one_hot_167709[27], one_hot_167709[1] | one_hot_167709[3] | one_hot_167709[5] | one_hot_167709[7] | one_hot_167709[9] | one_hot_167709[11] | one_hot_167709[13] | one_hot_167709[15] | one_hot_167709[17] | one_hot_167709[19] | one_hot_167709[21] | one_hot_167709[23] | one_hot_167709[25] | one_hot_167709[27]};
  assign one_hot_167718 = {reverse_167710[27:0] == 28'h000_0000, reverse_167710[27] && reverse_167710[26:0] == 27'h000_0000, reverse_167710[26] && reverse_167710[25:0] == 26'h000_0000, reverse_167710[25] && reverse_167710[24:0] == 25'h000_0000, reverse_167710[24] && reverse_167710[23:0] == 24'h00_0000, reverse_167710[23] && reverse_167710[22:0] == 23'h00_0000, reverse_167710[22] && reverse_167710[21:0] == 22'h00_0000, reverse_167710[21] && reverse_167710[20:0] == 21'h00_0000, reverse_167710[20] && reverse_167710[19:0] == 20'h0_0000, reverse_167710[19] && reverse_167710[18:0] == 19'h0_0000, reverse_167710[18] && reverse_167710[17:0] == 18'h0_0000, reverse_167710[17] && reverse_167710[16:0] == 17'h0_0000, reverse_167710[16] && reverse_167710[15:0] == 16'h0000, reverse_167710[15] && reverse_167710[14:0] == 15'h0000, reverse_167710[14] && reverse_167710[13:0] == 14'h0000, reverse_167710[13] && reverse_167710[12:0] == 13'h0000, reverse_167710[12] && reverse_167710[11:0] == 12'h000, reverse_167710[11] && reverse_167710[10:0] == 11'h000, reverse_167710[10] && reverse_167710[9:0] == 10'h000, reverse_167710[9] && reverse_167710[8:0] == 9'h000, reverse_167710[8] && reverse_167710[7:0] == 8'h00, reverse_167710[7] && reverse_167710[6:0] == 7'h00, reverse_167710[6] && reverse_167710[5:0] == 6'h00, reverse_167710[5] && reverse_167710[4:0] == 5'h00, reverse_167710[4] && reverse_167710[3:0] == 4'h0, reverse_167710[3] && reverse_167710[2:0] == 3'h0, reverse_167710[2] && reverse_167710[1:0] == 2'h0, reverse_167710[1] && !reverse_167710[0], reverse_167710[0]};
  assign encode_167719 = {one_hot_167711[16] | one_hot_167711[17] | one_hot_167711[18] | one_hot_167711[19] | one_hot_167711[20] | one_hot_167711[21] | one_hot_167711[22] | one_hot_167711[23] | one_hot_167711[24] | one_hot_167711[25] | one_hot_167711[26] | one_hot_167711[27] | one_hot_167711[28], one_hot_167711[8] | one_hot_167711[9] | one_hot_167711[10] | one_hot_167711[11] | one_hot_167711[12] | one_hot_167711[13] | one_hot_167711[14] | one_hot_167711[15] | one_hot_167711[24] | one_hot_167711[25] | one_hot_167711[26] | one_hot_167711[27] | one_hot_167711[28], one_hot_167711[4] | one_hot_167711[5] | one_hot_167711[6] | one_hot_167711[7] | one_hot_167711[12] | one_hot_167711[13] | one_hot_167711[14] | one_hot_167711[15] | one_hot_167711[20] | one_hot_167711[21] | one_hot_167711[22] | one_hot_167711[23] | one_hot_167711[28], one_hot_167711[2] | one_hot_167711[3] | one_hot_167711[6] | one_hot_167711[7] | one_hot_167711[10] | one_hot_167711[11] | one_hot_167711[14] | one_hot_167711[15] | one_hot_167711[18] | one_hot_167711[19] | one_hot_167711[22] | one_hot_167711[23] | one_hot_167711[26] | one_hot_167711[27], one_hot_167711[1] | one_hot_167711[3] | one_hot_167711[5] | one_hot_167711[7] | one_hot_167711[9] | one_hot_167711[11] | one_hot_167711[13] | one_hot_167711[15] | one_hot_167711[17] | one_hot_167711[19] | one_hot_167711[21] | one_hot_167711[23] | one_hot_167711[25] | one_hot_167711[27]};
  assign one_hot_167720 = {reverse_167712[27:0] == 28'h000_0000, reverse_167712[27] && reverse_167712[26:0] == 27'h000_0000, reverse_167712[26] && reverse_167712[25:0] == 26'h000_0000, reverse_167712[25] && reverse_167712[24:0] == 25'h000_0000, reverse_167712[24] && reverse_167712[23:0] == 24'h00_0000, reverse_167712[23] && reverse_167712[22:0] == 23'h00_0000, reverse_167712[22] && reverse_167712[21:0] == 22'h00_0000, reverse_167712[21] && reverse_167712[20:0] == 21'h00_0000, reverse_167712[20] && reverse_167712[19:0] == 20'h0_0000, reverse_167712[19] && reverse_167712[18:0] == 19'h0_0000, reverse_167712[18] && reverse_167712[17:0] == 18'h0_0000, reverse_167712[17] && reverse_167712[16:0] == 17'h0_0000, reverse_167712[16] && reverse_167712[15:0] == 16'h0000, reverse_167712[15] && reverse_167712[14:0] == 15'h0000, reverse_167712[14] && reverse_167712[13:0] == 14'h0000, reverse_167712[13] && reverse_167712[12:0] == 13'h0000, reverse_167712[12] && reverse_167712[11:0] == 12'h000, reverse_167712[11] && reverse_167712[10:0] == 11'h000, reverse_167712[10] && reverse_167712[9:0] == 10'h000, reverse_167712[9] && reverse_167712[8:0] == 9'h000, reverse_167712[8] && reverse_167712[7:0] == 8'h00, reverse_167712[7] && reverse_167712[6:0] == 7'h00, reverse_167712[6] && reverse_167712[5:0] == 6'h00, reverse_167712[5] && reverse_167712[4:0] == 5'h00, reverse_167712[4] && reverse_167712[3:0] == 4'h0, reverse_167712[3] && reverse_167712[2:0] == 3'h0, reverse_167712[2] && reverse_167712[1:0] == 2'h0, reverse_167712[1] && !reverse_167712[0], reverse_167712[0]};
  assign encode_167721 = {one_hot_167713[16] | one_hot_167713[17] | one_hot_167713[18] | one_hot_167713[19] | one_hot_167713[20] | one_hot_167713[21] | one_hot_167713[22] | one_hot_167713[23] | one_hot_167713[24] | one_hot_167713[25] | one_hot_167713[26] | one_hot_167713[27] | one_hot_167713[28], one_hot_167713[8] | one_hot_167713[9] | one_hot_167713[10] | one_hot_167713[11] | one_hot_167713[12] | one_hot_167713[13] | one_hot_167713[14] | one_hot_167713[15] | one_hot_167713[24] | one_hot_167713[25] | one_hot_167713[26] | one_hot_167713[27] | one_hot_167713[28], one_hot_167713[4] | one_hot_167713[5] | one_hot_167713[6] | one_hot_167713[7] | one_hot_167713[12] | one_hot_167713[13] | one_hot_167713[14] | one_hot_167713[15] | one_hot_167713[20] | one_hot_167713[21] | one_hot_167713[22] | one_hot_167713[23] | one_hot_167713[28], one_hot_167713[2] | one_hot_167713[3] | one_hot_167713[6] | one_hot_167713[7] | one_hot_167713[10] | one_hot_167713[11] | one_hot_167713[14] | one_hot_167713[15] | one_hot_167713[18] | one_hot_167713[19] | one_hot_167713[22] | one_hot_167713[23] | one_hot_167713[26] | one_hot_167713[27], one_hot_167713[1] | one_hot_167713[3] | one_hot_167713[5] | one_hot_167713[7] | one_hot_167713[9] | one_hot_167713[11] | one_hot_167713[13] | one_hot_167713[15] | one_hot_167713[17] | one_hot_167713[19] | one_hot_167713[21] | one_hot_167713[23] | one_hot_167713[25] | one_hot_167713[27]};
  assign encode_167722 = {one_hot_167714[16] | one_hot_167714[17] | one_hot_167714[18] | one_hot_167714[19] | one_hot_167714[20] | one_hot_167714[21] | one_hot_167714[22] | one_hot_167714[23] | one_hot_167714[24] | one_hot_167714[25] | one_hot_167714[26] | one_hot_167714[27] | one_hot_167714[28], one_hot_167714[8] | one_hot_167714[9] | one_hot_167714[10] | one_hot_167714[11] | one_hot_167714[12] | one_hot_167714[13] | one_hot_167714[14] | one_hot_167714[15] | one_hot_167714[24] | one_hot_167714[25] | one_hot_167714[26] | one_hot_167714[27] | one_hot_167714[28], one_hot_167714[4] | one_hot_167714[5] | one_hot_167714[6] | one_hot_167714[7] | one_hot_167714[12] | one_hot_167714[13] | one_hot_167714[14] | one_hot_167714[15] | one_hot_167714[20] | one_hot_167714[21] | one_hot_167714[22] | one_hot_167714[23] | one_hot_167714[28], one_hot_167714[2] | one_hot_167714[3] | one_hot_167714[6] | one_hot_167714[7] | one_hot_167714[10] | one_hot_167714[11] | one_hot_167714[14] | one_hot_167714[15] | one_hot_167714[18] | one_hot_167714[19] | one_hot_167714[22] | one_hot_167714[23] | one_hot_167714[26] | one_hot_167714[27], one_hot_167714[1] | one_hot_167714[3] | one_hot_167714[5] | one_hot_167714[7] | one_hot_167714[9] | one_hot_167714[11] | one_hot_167714[13] | one_hot_167714[15] | one_hot_167714[17] | one_hot_167714[19] | one_hot_167714[21] | one_hot_167714[23] | one_hot_167714[25] | one_hot_167714[27]};
  assign encode_167724 = {one_hot_167716[16] | one_hot_167716[17] | one_hot_167716[18] | one_hot_167716[19] | one_hot_167716[20] | one_hot_167716[21] | one_hot_167716[22] | one_hot_167716[23] | one_hot_167716[24] | one_hot_167716[25] | one_hot_167716[26] | one_hot_167716[27] | one_hot_167716[28], one_hot_167716[8] | one_hot_167716[9] | one_hot_167716[10] | one_hot_167716[11] | one_hot_167716[12] | one_hot_167716[13] | one_hot_167716[14] | one_hot_167716[15] | one_hot_167716[24] | one_hot_167716[25] | one_hot_167716[26] | one_hot_167716[27] | one_hot_167716[28], one_hot_167716[4] | one_hot_167716[5] | one_hot_167716[6] | one_hot_167716[7] | one_hot_167716[12] | one_hot_167716[13] | one_hot_167716[14] | one_hot_167716[15] | one_hot_167716[20] | one_hot_167716[21] | one_hot_167716[22] | one_hot_167716[23] | one_hot_167716[28], one_hot_167716[2] | one_hot_167716[3] | one_hot_167716[6] | one_hot_167716[7] | one_hot_167716[10] | one_hot_167716[11] | one_hot_167716[14] | one_hot_167716[15] | one_hot_167716[18] | one_hot_167716[19] | one_hot_167716[22] | one_hot_167716[23] | one_hot_167716[26] | one_hot_167716[27], one_hot_167716[1] | one_hot_167716[3] | one_hot_167716[5] | one_hot_167716[7] | one_hot_167716[9] | one_hot_167716[11] | one_hot_167716[13] | one_hot_167716[15] | one_hot_167716[17] | one_hot_167716[19] | one_hot_167716[21] | one_hot_167716[23] | one_hot_167716[25] | one_hot_167716[27]};
  assign encode_167726 = {one_hot_167718[16] | one_hot_167718[17] | one_hot_167718[18] | one_hot_167718[19] | one_hot_167718[20] | one_hot_167718[21] | one_hot_167718[22] | one_hot_167718[23] | one_hot_167718[24] | one_hot_167718[25] | one_hot_167718[26] | one_hot_167718[27] | one_hot_167718[28], one_hot_167718[8] | one_hot_167718[9] | one_hot_167718[10] | one_hot_167718[11] | one_hot_167718[12] | one_hot_167718[13] | one_hot_167718[14] | one_hot_167718[15] | one_hot_167718[24] | one_hot_167718[25] | one_hot_167718[26] | one_hot_167718[27] | one_hot_167718[28], one_hot_167718[4] | one_hot_167718[5] | one_hot_167718[6] | one_hot_167718[7] | one_hot_167718[12] | one_hot_167718[13] | one_hot_167718[14] | one_hot_167718[15] | one_hot_167718[20] | one_hot_167718[21] | one_hot_167718[22] | one_hot_167718[23] | one_hot_167718[28], one_hot_167718[2] | one_hot_167718[3] | one_hot_167718[6] | one_hot_167718[7] | one_hot_167718[10] | one_hot_167718[11] | one_hot_167718[14] | one_hot_167718[15] | one_hot_167718[18] | one_hot_167718[19] | one_hot_167718[22] | one_hot_167718[23] | one_hot_167718[26] | one_hot_167718[27], one_hot_167718[1] | one_hot_167718[3] | one_hot_167718[5] | one_hot_167718[7] | one_hot_167718[9] | one_hot_167718[11] | one_hot_167718[13] | one_hot_167718[15] | one_hot_167718[17] | one_hot_167718[19] | one_hot_167718[21] | one_hot_167718[23] | one_hot_167718[25] | one_hot_167718[27]};
  assign encode_167728 = {one_hot_167720[16] | one_hot_167720[17] | one_hot_167720[18] | one_hot_167720[19] | one_hot_167720[20] | one_hot_167720[21] | one_hot_167720[22] | one_hot_167720[23] | one_hot_167720[24] | one_hot_167720[25] | one_hot_167720[26] | one_hot_167720[27] | one_hot_167720[28], one_hot_167720[8] | one_hot_167720[9] | one_hot_167720[10] | one_hot_167720[11] | one_hot_167720[12] | one_hot_167720[13] | one_hot_167720[14] | one_hot_167720[15] | one_hot_167720[24] | one_hot_167720[25] | one_hot_167720[26] | one_hot_167720[27] | one_hot_167720[28], one_hot_167720[4] | one_hot_167720[5] | one_hot_167720[6] | one_hot_167720[7] | one_hot_167720[12] | one_hot_167720[13] | one_hot_167720[14] | one_hot_167720[15] | one_hot_167720[20] | one_hot_167720[21] | one_hot_167720[22] | one_hot_167720[23] | one_hot_167720[28], one_hot_167720[2] | one_hot_167720[3] | one_hot_167720[6] | one_hot_167720[7] | one_hot_167720[10] | one_hot_167720[11] | one_hot_167720[14] | one_hot_167720[15] | one_hot_167720[18] | one_hot_167720[19] | one_hot_167720[22] | one_hot_167720[23] | one_hot_167720[26] | one_hot_167720[27], one_hot_167720[1] | one_hot_167720[3] | one_hot_167720[5] | one_hot_167720[7] | one_hot_167720[9] | one_hot_167720[11] | one_hot_167720[13] | one_hot_167720[15] | one_hot_167720[17] | one_hot_167720[19] | one_hot_167720[21] | one_hot_167720[23] | one_hot_167720[25] | one_hot_167720[27]};
  assign cancel__16 = |encode_167715[4:1];
  assign carry_bit__15 = xbs_fraction__15[27];
  assign result_fraction__514 = 23'h00_0000;
  assign cancel__32 = |encode_167717[4:1];
  assign carry_bit__32 = xbs_fraction__31[27];
  assign result_fraction__581 = 23'h00_0000;
  assign cancel__51 = |encode_167719[4:1];
  assign carry_bit__51 = xbs_fraction__49[27];
  assign result_fraction__648 = 23'h00_0000;
  assign cancel__70 = |encode_167721[4:1];
  assign carry_bit__70 = xbs_fraction__67[27];
  assign result_fraction__723 = 23'h00_0000;
  assign cancel__7 = |encode_167722[4:1];
  assign carry_bit__7 = xbs_fraction__7[27];
  assign result_fraction__515 = 23'h00_0000;
  assign leading_zeroes__15 = {result_fraction__514, encode_167715};
  assign cancel__33 = |encode_167724[4:1];
  assign carry_bit__33 = xbs_fraction__32[27];
  assign result_fraction__582 = 23'h00_0000;
  assign leading_zeroes__32 = {result_fraction__581, encode_167717};
  assign cancel__52 = |encode_167726[4:1];
  assign carry_bit__52 = xbs_fraction__50[27];
  assign result_fraction__649 = 23'h00_0000;
  assign leading_zeroes__51 = {result_fraction__648, encode_167719};
  assign cancel__71 = |encode_167728[4:1];
  assign carry_bit__71 = xbs_fraction__68[27];
  assign result_fraction__724 = 23'h00_0000;
  assign leading_zeroes__70 = {result_fraction__723, encode_167721};
  assign array_index_167783 = in_img_unflattened[4'he];
  assign leading_zeroes__7 = {result_fraction__515, encode_167722};
  assign carry_fraction__30 = xbs_fraction__15[27:1];
  assign add_167796 = leading_zeroes__15 + 28'hfff_ffff;
  assign leading_zeroes__33 = {result_fraction__582, encode_167724};
  assign carry_fraction__63 = xbs_fraction__31[27:1];
  assign add_167809 = leading_zeroes__32 + 28'hfff_ffff;
  assign leading_zeroes__52 = {result_fraction__649, encode_167726};
  assign carry_fraction__101 = xbs_fraction__49[27:1];
  assign add_167822 = leading_zeroes__51 + 28'hfff_ffff;
  assign leading_zeroes__71 = {result_fraction__724, encode_167728};
  assign carry_fraction__139 = xbs_fraction__67[27:1];
  assign add_167835 = leading_zeroes__70 + 28'hfff_ffff;
  assign x_bexp__541 = array_index_167783[30:23];
  assign carry_fraction__13 = xbs_fraction__7[27:1];
  assign add_167843 = leading_zeroes__7 + 28'hfff_ffff;
  assign concat_167844 = {~(carry_bit__15 | cancel__16), ~(carry_bit__15 | ~cancel__16), ~(~carry_bit__15 | cancel__16)};
  assign carry_fraction__31 = carry_fraction__30 | {26'h000_0000, xbs_fraction__15[0]};
  assign cancel_fraction__15 = add_167796 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__15[26:0] << add_167796;
  assign carry_fraction__64 = xbs_fraction__32[27:1];
  assign add_167853 = leading_zeroes__33 + 28'hfff_ffff;
  assign concat_167854 = {~(carry_bit__32 | cancel__32), ~(carry_bit__32 | ~cancel__32), ~(~carry_bit__32 | cancel__32)};
  assign carry_fraction__65 = carry_fraction__63 | {26'h000_0000, xbs_fraction__31[0]};
  assign cancel_fraction__32 = add_167809 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__31[26:0] << add_167809;
  assign carry_fraction__102 = xbs_fraction__50[27:1];
  assign add_167863 = leading_zeroes__52 + 28'hfff_ffff;
  assign concat_167864 = {~(carry_bit__51 | cancel__51), ~(carry_bit__51 | ~cancel__51), ~(~carry_bit__51 | cancel__51)};
  assign carry_fraction__103 = carry_fraction__101 | {26'h000_0000, xbs_fraction__49[0]};
  assign cancel_fraction__51 = add_167822 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__49[26:0] << add_167822;
  assign result_sign__1058 = 1'h0;
  assign carry_fraction__140 = xbs_fraction__68[27:1];
  assign add_167875 = leading_zeroes__71 + 28'hfff_ffff;
  assign concat_167876 = {~(carry_bit__70 | cancel__70), ~(carry_bit__70 | ~cancel__70), ~(~carry_bit__70 | cancel__70)};
  assign carry_fraction__141 = carry_fraction__139 | {26'h000_0000, xbs_fraction__67[0]};
  assign cancel_fraction__70 = add_167835 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__67[26:0] << add_167835;
  assign result_sign__1059 = 1'h0;
  assign concat_167881 = {~(carry_bit__7 | cancel__7), ~(carry_bit__7 | ~cancel__7), ~(~carry_bit__7 | cancel__7)};
  assign carry_fraction__14 = carry_fraction__13 | {26'h000_0000, xbs_fraction__7[0]};
  assign cancel_fraction__7 = add_167843 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__7[26:0] << add_167843;
  assign shifted_fraction__15 = carry_fraction__31 & {27{concat_167844[0]}} | cancel_fraction__15 & {27{concat_167844[1]}} | xbs_fraction__15[26:0] & {27{concat_167844[2]}};
  assign concat_167885 = {~(carry_bit__33 | cancel__33), ~(carry_bit__33 | ~cancel__33), ~(~carry_bit__33 | cancel__33)};
  assign carry_fraction__66 = carry_fraction__64 | {26'h000_0000, xbs_fraction__32[0]};
  assign cancel_fraction__33 = add_167853 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__32[26:0] << add_167853;
  assign shifted_fraction__32 = carry_fraction__65 & {27{concat_167854[0]}} | cancel_fraction__32 & {27{concat_167854[1]}} | xbs_fraction__31[26:0] & {27{concat_167854[2]}};
  assign concat_167889 = {~(carry_bit__52 | cancel__52), ~(carry_bit__52 | ~cancel__52), ~(~carry_bit__52 | cancel__52)};
  assign carry_fraction__104 = carry_fraction__102 | {26'h000_0000, xbs_fraction__50[0]};
  assign cancel_fraction__52 = add_167863 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__50[26:0] << add_167863;
  assign shifted_fraction__51 = carry_fraction__103 & {27{concat_167864[0]}} | cancel_fraction__51 & {27{concat_167864[1]}} | xbs_fraction__49[26:0] & {27{concat_167864[2]}};
  assign concat_167895 = {~(carry_bit__71 | cancel__71), ~(carry_bit__71 | ~cancel__71), ~(~carry_bit__71 | cancel__71)};
  assign carry_fraction__142 = carry_fraction__140 | {26'h000_0000, xbs_fraction__68[0]};
  assign cancel_fraction__71 = add_167875 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__68[26:0] << add_167875;
  assign shifted_fraction__70 = carry_fraction__141 & {27{concat_167876[0]}} | cancel_fraction__70 & {27{concat_167876[1]}} | xbs_fraction__67[26:0] & {27{concat_167876[2]}};
  assign shifted_fraction__7 = carry_fraction__14 & {27{concat_167881[0]}} | cancel_fraction__7 & {27{concat_167881[1]}} | xbs_fraction__7[26:0] & {27{concat_167881[2]}};
  assign result_sign__1060 = 1'h0;
  assign shifted_fraction__33 = carry_fraction__66 & {27{concat_167885[0]}} | cancel_fraction__33 & {27{concat_167885[1]}} | xbs_fraction__32[26:0] & {27{concat_167885[2]}};
  assign result_sign__1061 = 1'h0;
  assign shifted_fraction__52 = carry_fraction__104 & {27{concat_167889[0]}} | cancel_fraction__52 & {27{concat_167889[1]}} | xbs_fraction__50[26:0] & {27{concat_167889[2]}};
  assign result_sign__1062 = 1'h0;
  assign result_sign__1111 = 1'h0;
  assign add_167911 = {result_sign__1058, x_bexp__525[7]} + 2'h1;
  assign shifted_fraction__71 = carry_fraction__142 & {27{concat_167895[0]}} | cancel_fraction__71 & {27{concat_167895[1]}} | xbs_fraction__68[26:0] & {27{concat_167895[2]}};
  assign result_sign__1063 = 1'h0;
  assign result_sign__1115 = 1'h0;
  assign add_167917 = {result_sign__1059, x_bexp__541[7]} + 2'h1;
  assign x_bexp__778 = 8'h00;
  assign result_sign__747 = 1'h0;
  assign x_fraction__541 = array_index_167783[22:0];
  assign result_sign__1064 = 1'h0;
  assign normal_chunk__15 = shifted_fraction__15[2:0];
  assign fraction_shift__249 = 3'h4;
  assign half_way_chunk__15 = shifted_fraction__15[3:2];
  assign result_sign__1065 = 1'h0;
  assign normal_chunk__32 = shifted_fraction__32[2:0];
  assign fraction_shift__284 = 3'h4;
  assign half_way_chunk__32 = shifted_fraction__32[3:2];
  assign result_sign__1066 = 1'h0;
  assign normal_chunk__51 = shifted_fraction__51[2:0];
  assign fraction_shift__319 = 3'h4;
  assign half_way_chunk__51 = shifted_fraction__51[3:2];
  assign result_sign__1067 = 1'h0;
  assign normal_chunk__70 = shifted_fraction__70[2:0];
  assign fraction_shift__354 = 3'h4;
  assign half_way_chunk__70 = shifted_fraction__70[3:2];
  assign ne_167958 = x_bexp__541 != x_bexp__778;
  assign normal_chunk__7 = shifted_fraction__7[2:0];
  assign fraction_shift__250 = 3'h4;
  assign half_way_chunk__7 = shifted_fraction__7[3:2];
  assign result_sign__442 = 1'h0;
  assign add_167970 = {result_sign__1060, shifted_fraction__15[26:3]} + 25'h000_0001;
  assign normal_chunk__33 = shifted_fraction__33[2:0];
  assign fraction_shift__285 = 3'h4;
  assign half_way_chunk__33 = shifted_fraction__33[3:2];
  assign result_sign__539 = 1'h0;
  assign add_167980 = {result_sign__1061, shifted_fraction__32[26:3]} + 25'h000_0001;
  assign normal_chunk__52 = shifted_fraction__52[2:0];
  assign fraction_shift__320 = 3'h4;
  assign half_way_chunk__52 = shifted_fraction__52[3:2];
  assign result_sign__639 = 1'h0;
  assign add_167990 = {result_sign__1062, shifted_fraction__51[26:3]} + 25'h000_0001;
  assign exp__221 = {result_sign__1111, add_167911, x_bexp__525[6:0]} + 10'h381;
  assign normal_chunk__71 = shifted_fraction__71[2:0];
  assign fraction_shift__355 = 3'h4;
  assign half_way_chunk__71 = shifted_fraction__71[3:2];
  assign result_sign__749 = 1'h0;
  assign add_168001 = {result_sign__1063, shifted_fraction__70[26:3]} + 25'h000_0001;
  assign exp__303 = {result_sign__1115, add_167917, x_bexp__541[6:0]} + 10'h381;
  assign sign_ext_168003 = {10{ne_167958}};
  assign x_fraction__543 = {result_sign__747, x_fraction__541} | 24'h80_0000;
  assign result_sign__443 = 1'h0;
  assign add_168009 = {result_sign__1064, shifted_fraction__7[26:3]} + 25'h000_0001;
  assign do_round_up__31 = normal_chunk__15 > fraction_shift__249 | half_way_chunk__15 == 2'h3;
  assign result_sign__540 = 1'h0;
  assign add_168016 = {result_sign__1065, shifted_fraction__33[26:3]} + 25'h000_0001;
  assign do_round_up__66 = normal_chunk__32 > fraction_shift__284 | half_way_chunk__32 == 2'h3;
  assign result_sign__640 = 1'h0;
  assign add_168023 = {result_sign__1066, shifted_fraction__52[26:3]} + 25'h000_0001;
  assign do_round_up__105 = normal_chunk__51 > fraction_shift__319 | half_way_chunk__51 == 2'h3;
  assign exp__223 = exp__221 & sign_ext_166301;
  assign result_sign__750 = 1'h0;
  assign add_168032 = {result_sign__1067, shifted_fraction__71[26:3]} + 25'h000_0001;
  assign do_round_up__144 = normal_chunk__70 > fraction_shift__354 | half_way_chunk__70 == 2'h3;
  assign exp__305 = exp__303 & sign_ext_168003;
  assign x_fraction__545 = x_fraction__543 & {24{ne_167958}};
  assign result_sign__824 = 1'h0;
  assign result_sign__825 = 1'h0;
  assign do_round_up__14 = normal_chunk__7 > fraction_shift__250 | half_way_chunk__7 == 2'h3;
  assign rounded_fraction__15 = do_round_up__31 ? {add_167970, normal_chunk__15} : {result_sign__442, shifted_fraction__15};
  assign do_round_up__67 = normal_chunk__33 > fraction_shift__285 | half_way_chunk__33 == 2'h3;
  assign rounded_fraction__32 = do_round_up__66 ? {add_167980, normal_chunk__32} : {result_sign__539, shifted_fraction__32};
  assign do_round_up__106 = normal_chunk__52 > fraction_shift__320 | half_way_chunk__52 == 2'h3;
  assign rounded_fraction__51 = do_round_up__105 ? {add_167990, normal_chunk__51} : {result_sign__639, shifted_fraction__51};
  assign do_round_up__145 = normal_chunk__71 > fraction_shift__355 | half_way_chunk__71 == 2'h3;
  assign rounded_fraction__70 = do_round_up__144 ? {add_168001, normal_chunk__70} : {result_sign__749, shifted_fraction__70};
  assign concat_168059 = {x_fraction__545, result_sign__824};
  assign concat_168060 = {result_sign__825, x_fraction__545};
  assign rounded_fraction__7 = do_round_up__14 ? {add_168009, normal_chunk__7} : {result_sign__443, shifted_fraction__7};
  assign result_sign__444 = 1'h0;
  assign x_bexp__586 = 8'h00;
  assign rounding_carry__15 = rounded_fraction__15[27];
  assign rounded_fraction__33 = do_round_up__67 ? {add_168016, normal_chunk__33} : {result_sign__540, shifted_fraction__33};
  assign result_sign__541 = 1'h0;
  assign x_bexp__604 = 8'h00;
  assign rounding_carry__32 = rounded_fraction__32[27];
  assign rounded_fraction__52 = do_round_up__106 ? {add_168023, normal_chunk__52} : {result_sign__640, shifted_fraction__52};
  assign result_sign__641 = 1'h0;
  assign x_bexp__622 = 8'h00;
  assign rounding_carry__51 = rounded_fraction__51[27];
  assign sel_168073 = $signed(exp__223) <= $signed(10'h000) ? concat_166369 : concat_166368;
  assign rounded_fraction__71 = do_round_up__145 ? {add_168032, normal_chunk__71} : {result_sign__750, shifted_fraction__71};
  assign result_sign__751 = 1'h0;
  assign x_bexp__640 = 8'h00;
  assign rounding_carry__70 = rounded_fraction__70[27];
  assign sel_168078 = $signed(exp__305) <= $signed(10'h000) ? concat_168060 : concat_168059;
  assign result_sign__445 = 1'h0;
  assign x_bexp__587 = 8'h00;
  assign rounding_carry__7 = rounded_fraction__7[27];
  assign result_sign__542 = 1'h0;
  assign x_bexp__605 = 8'h00;
  assign rounding_carry__33 = rounded_fraction__33[27];
  assign result_sign__642 = 1'h0;
  assign x_bexp__623 = 8'h00;
  assign rounding_carry__52 = rounded_fraction__52[27];
  assign result_sign__946 = 1'h0;
  assign fraction__495 = sel_168073[23:1];
  assign result_sign__752 = 1'h0;
  assign x_bexp__641 = 8'h00;
  assign rounding_carry__71 = rounded_fraction__71[27];
  assign result_sign__954 = 1'h0;
  assign fraction__674 = sel_168078[23:1];
  assign result_sign__446 = 1'h0;
  assign add_168106 = {result_sign__444, x_bexp__126} + {x_bexp__586, rounding_carry__15};
  assign result_sign__543 = 1'h0;
  assign add_168112 = {result_sign__541, x_bexp__251} + {x_bexp__604, rounding_carry__32};
  assign result_sign__643 = 1'h0;
  assign add_168118 = {result_sign__641, x_bexp__395} + {x_bexp__622, rounding_carry__51};
  assign fraction__497 = {result_sign__946, fraction__495};
  assign result_sign__753 = 1'h0;
  assign add_168128 = {result_sign__751, x_bexp__539} + {x_bexp__640, rounding_carry__70};
  assign fraction__676 = {result_sign__954, fraction__674};
  assign result_sign__447 = 1'h0;
  assign add_168136 = {result_sign__445, x_bexp__54} + {x_bexp__587, rounding_carry__7};
  assign result_sign__544 = 1'h0;
  assign add_168145 = {result_sign__542, x_bexp__252} + {x_bexp__605, rounding_carry__33};
  assign result_sign__644 = 1'h0;
  assign add_168154 = {result_sign__642, x_bexp__396} + {x_bexp__623, rounding_carry__52};
  assign do_round_up__107 = sel_168073[0] & sel_168073[1];
  assign add_168163 = fraction__497 + 24'h00_0001;
  assign result_sign__754 = 1'h0;
  assign add_168165 = {result_sign__752, x_bexp__540} + {x_bexp__641, rounding_carry__71};
  assign do_round_up__146 = sel_168078[0] & sel_168078[1];
  assign add_168174 = fraction__676 + 24'h00_0001;
  assign add_168180 = {result_sign__446, add_168106} + 10'h001;
  assign add_168188 = {result_sign__543, add_168112} + 10'h001;
  assign add_168196 = {result_sign__643, add_168118} + 10'h001;
  assign fraction__499 = do_round_up__107 ? add_168163 : fraction__497;
  assign add_168206 = {result_sign__753, add_168128} + 10'h001;
  assign fraction__678 = do_round_up__146 ? add_168174 : fraction__676;
  assign add_168211 = {result_sign__447, add_168136} + 10'h001;
  assign wide_exponent__45 = add_168180 - {5'h00, encode_167715};
  assign add_168216 = {result_sign__544, add_168145} + 10'h001;
  assign wide_exponent__94 = add_168188 - {5'h00, encode_167717};
  assign add_168221 = {result_sign__644, add_168154} + 10'h001;
  assign wide_exponent__151 = add_168196 - {5'h00, encode_167719};
  assign add_168227 = exp__223 + 10'h001;
  assign add_168228 = {result_sign__754, add_168165} + 10'h001;
  assign wide_exponent__208 = add_168206 - {5'h00, encode_167721};
  assign add_168234 = exp__305 + 10'h001;
  assign wide_exponent__19 = add_168211 - {5'h00, encode_167722};
  assign wide_exponent__46 = wide_exponent__45 & {10{add_167640 != 26'h000_0000 | xddend_y__15[2:0] != 3'h0}};
  assign wide_exponent__95 = add_168216 - {5'h00, encode_167724};
  assign wide_exponent__96 = wide_exponent__94 & {10{add_167643 != 26'h000_0000 | xddend_y__31[2:0] != 3'h0}};
  assign wide_exponent__152 = add_168221 - {5'h00, encode_167726};
  assign wide_exponent__153 = wide_exponent__151 & {10{add_167646 != 26'h000_0000 | xddend_y__49[2:0] != 3'h0}};
  assign exp__227 = fraction__499[23] ? add_168227 : exp__223;
  assign wide_exponent__209 = add_168228 - {5'h00, encode_167728};
  assign wide_exponent__210 = wide_exponent__208 & {10{add_167649 != 26'h000_0000 | xddend_y__67[2:0] != 3'h0}};
  assign exp__309 = fraction__678[23] ? add_168234 : exp__305;
  assign wide_exponent__20 = wide_exponent__19 & {10{add_167650 != 26'h000_0000 | xddend_y__7[2:0] != 3'h0}};
  assign high_exp__375 = 8'hff;
  assign result_fraction__781 = 23'h00_0000;
  assign high_exp__376 = 8'hff;
  assign result_fraction__782 = 23'h00_0000;
  assign high_exp__117 = 8'hff;
  assign result_fraction__516 = 23'h00_0000;
  assign high_exp__118 = 8'hff;
  assign result_fraction__517 = 23'h00_0000;
  assign wide_exponent__97 = wide_exponent__95 & {10{add_167653 != 26'h000_0000 | xddend_y__32[2:0] != 3'h0}};
  assign high_exp__407 = 8'hff;
  assign result_fraction__814 = 23'h00_0000;
  assign high_exp__408 = 8'hff;
  assign result_fraction__815 = 23'h00_0000;
  assign high_exp__182 = 8'hff;
  assign result_fraction__583 = 23'h00_0000;
  assign high_exp__183 = 8'hff;
  assign result_fraction__584 = 23'h00_0000;
  assign wide_exponent__154 = wide_exponent__152 & {10{add_167656 != 26'h000_0000 | xddend_y__50[2:0] != 3'h0}};
  assign high_exp__439 = 8'hff;
  assign result_fraction__847 = 23'h00_0000;
  assign high_exp__440 = 8'hff;
  assign result_fraction__848 = 23'h00_0000;
  assign high_exp__249 = 8'hff;
  assign result_fraction__650 = 23'h00_0000;
  assign high_exp__250 = 8'hff;
  assign result_fraction__651 = 23'h00_0000;
  assign wide_exponent__211 = wide_exponent__209 & {10{add_167659 != 26'h000_0000 | xddend_y__68[2:0] != 3'h0}};
  assign high_exp__471 = 8'hff;
  assign result_fraction__880 = 23'h00_0000;
  assign high_exp__472 = 8'hff;
  assign result_fraction__881 = 23'h00_0000;
  assign high_exp__321 = 8'hff;
  assign result_fraction__725 = 23'h00_0000;
  assign high_exp__322 = 8'hff;
  assign result_fraction__726 = 23'h00_0000;
  assign high_exp__361 = 8'hff;
  assign result_fraction__766 = 23'h00_0000;
  assign high_exp__362 = 8'hff;
  assign result_fraction__767 = 23'h00_0000;
  assign high_exp__119 = 8'hff;
  assign result_fraction__518 = 23'h00_0000;
  assign high_exp__120 = 8'hff;
  assign result_fraction__519 = 23'h00_0000;
  assign ne_168304 = x_fraction__126 != result_fraction__781;
  assign ne_168306 = prod_fraction__45 != result_fraction__782;
  assign eq_168307 = x_bexp__126 == high_exp__117;
  assign eq_168308 = x_fraction__126 == result_fraction__516;
  assign eq_168309 = prod_bexp__62 == high_exp__118;
  assign eq_168310 = prod_fraction__45 == result_fraction__517;
  assign high_exp__393 = 8'hff;
  assign result_fraction__799 = 23'h00_0000;
  assign high_exp__394 = 8'hff;
  assign result_fraction__800 = 23'h00_0000;
  assign high_exp__184 = 8'hff;
  assign result_fraction__585 = 23'h00_0000;
  assign high_exp__185 = 8'hff;
  assign result_fraction__586 = 23'h00_0000;
  assign ne_168322 = x_fraction__251 != result_fraction__814;
  assign ne_168324 = prod_fraction__91 != result_fraction__815;
  assign eq_168325 = x_bexp__251 == high_exp__182;
  assign eq_168326 = x_fraction__251 == result_fraction__583;
  assign eq_168327 = prod_bexp__123 == high_exp__183;
  assign eq_168328 = prod_fraction__91 == result_fraction__584;
  assign high_exp__425 = 8'hff;
  assign result_fraction__832 = 23'h00_0000;
  assign high_exp__426 = 8'hff;
  assign result_fraction__833 = 23'h00_0000;
  assign high_exp__251 = 8'hff;
  assign result_fraction__652 = 23'h00_0000;
  assign high_exp__252 = 8'hff;
  assign result_fraction__653 = 23'h00_0000;
  assign ne_168340 = x_fraction__395 != result_fraction__847;
  assign ne_168342 = prod_fraction__145 != result_fraction__848;
  assign eq_168343 = x_bexp__395 == high_exp__249;
  assign eq_168344 = x_fraction__395 == result_fraction__650;
  assign eq_168345 = prod_bexp__195 == high_exp__250;
  assign eq_168346 = prod_fraction__145 == result_fraction__651;
  assign result_exp__163 = exp__227[8:0];
  assign high_exp__457 = 8'hff;
  assign result_fraction__865 = 23'h00_0000;
  assign high_exp__458 = 8'hff;
  assign result_fraction__866 = 23'h00_0000;
  assign high_exp__323 = 8'hff;
  assign result_fraction__727 = 23'h00_0000;
  assign high_exp__324 = 8'hff;
  assign result_fraction__728 = 23'h00_0000;
  assign ne_168360 = x_fraction__539 != result_fraction__880;
  assign ne_168362 = prod_fraction__199 != result_fraction__881;
  assign eq_168363 = x_bexp__539 == high_exp__321;
  assign eq_168364 = x_fraction__539 == result_fraction__725;
  assign eq_168365 = prod_bexp__267 == high_exp__322;
  assign eq_168366 = prod_fraction__199 == result_fraction__726;
  assign result_exp__223 = exp__309[8:0];
  assign ne_168371 = x_fraction__54 != result_fraction__766;
  assign ne_168373 = prod_fraction__19 != result_fraction__767;
  assign eq_168374 = x_bexp__54 == high_exp__119;
  assign eq_168375 = x_fraction__54 == result_fraction__518;
  assign eq_168376 = prod_bexp__26 == high_exp__120;
  assign eq_168377 = prod_fraction__19 == result_fraction__519;
  assign ne_168386 = x_fraction__252 != result_fraction__799;
  assign ne_168388 = prod_fraction__92 != result_fraction__800;
  assign eq_168389 = x_bexp__252 == high_exp__184;
  assign eq_168390 = x_fraction__252 == result_fraction__585;
  assign eq_168391 = prod_bexp__124 == high_exp__185;
  assign eq_168392 = prod_fraction__92 == result_fraction__586;
  assign ne_168401 = x_fraction__396 != result_fraction__832;
  assign ne_168403 = prod_fraction__146 != result_fraction__833;
  assign eq_168404 = x_bexp__396 == high_exp__251;
  assign eq_168405 = x_fraction__396 == result_fraction__652;
  assign eq_168406 = prod_bexp__196 == high_exp__252;
  assign eq_168407 = prod_fraction__146 == result_fraction__653;
  assign result_exp__165 = result_exp__163 & {9{$signed(exp__227) > $signed(10'h000)}};
  assign ne_168417 = x_fraction__540 != result_fraction__865;
  assign ne_168419 = prod_fraction__200 != result_fraction__866;
  assign eq_168420 = x_bexp__540 == high_exp__323;
  assign eq_168421 = x_fraction__540 == result_fraction__727;
  assign eq_168422 = prod_bexp__268 == high_exp__324;
  assign eq_168423 = prod_fraction__200 == result_fraction__728;
  assign high_exp__326 = 8'hff;
  assign result_fraction__730 = 23'h00_0000;
  assign result_fraction__729 = 23'h00_0000;
  assign result_exp__225 = result_exp__223 & {9{$signed(exp__309) > $signed(10'h000)}};
  assign wide_exponent__47 = wide_exponent__46[8:0] & {9{~wide_exponent__46[9]}};
  assign has_pos_inf__15 = ~(x_bexp__126 != high_exp__375 | ne_168304 | x_sign__32) | ~(prod_bexp__62 != high_exp__376 | ne_168306 | prod_sign__15);
  assign has_neg_inf__15 = eq_168307 & eq_168308 & x_sign__32 | eq_168309 & eq_168310 & prod_sign__15;
  assign wide_exponent__98 = wide_exponent__96[8:0] & {9{~wide_exponent__96[9]}};
  assign has_pos_inf__32 = ~(x_bexp__251 != high_exp__407 | ne_168322 | x_sign__63) | ~(prod_bexp__123 != high_exp__408 | ne_168324 | prod_sign__31);
  assign has_neg_inf__32 = eq_168325 & eq_168326 & x_sign__63 | eq_168327 & eq_168328 & prod_sign__31;
  assign wide_exponent__155 = wide_exponent__153[8:0] & {9{~wide_exponent__153[9]}};
  assign has_pos_inf__51 = ~(x_bexp__395 != high_exp__439 | ne_168340 | x_sign__99) | ~(prod_bexp__195 != high_exp__440 | ne_168342 | prod_sign__49);
  assign has_neg_inf__51 = eq_168343 & eq_168344 & x_sign__99 | eq_168345 & eq_168346 & prod_sign__49;
  assign wide_exponent__212 = wide_exponent__210[8:0] & {9{~wide_exponent__210[9]}};
  assign has_pos_inf__70 = ~(x_bexp__539 != high_exp__471 | ne_168360 | x_sign__135) | ~(prod_bexp__267 != high_exp__472 | ne_168362 | prod_sign__67);
  assign has_neg_inf__70 = eq_168363 & eq_168364 & x_sign__135 | eq_168365 & eq_168366 & prod_sign__67;
  assign is_result_nan__147 = x_bexp__541 == high_exp__326;
  assign ne_168472 = x_fraction__541 != result_fraction__730;
  assign wide_exponent__21 = wide_exponent__20[8:0] & {9{~wide_exponent__20[9]}};
  assign has_pos_inf__7 = ~(x_bexp__54 != high_exp__361 | ne_168371 | x_sign__14) | ~(prod_bexp__26 != high_exp__362 | ne_168373 | prod_sign__7);
  assign has_neg_inf__7 = eq_168374 & eq_168375 & x_sign__14 | eq_168376 & eq_168377 & prod_sign__7;
  assign wide_exponent__99 = wide_exponent__97[8:0] & {9{~wide_exponent__97[9]}};
  assign has_pos_inf__33 = ~(x_bexp__252 != high_exp__393 | ne_168386 | x_sign__64) | ~(prod_bexp__124 != high_exp__394 | ne_168388 | prod_sign__32);
  assign has_neg_inf__33 = eq_168389 & eq_168390 & x_sign__64 | eq_168391 & eq_168392 & prod_sign__32;
  assign wide_exponent__156 = wide_exponent__154[8:0] & {9{~wide_exponent__154[9]}};
  assign has_pos_inf__52 = ~(x_bexp__396 != high_exp__425 | ne_168401 | x_sign__100) | ~(prod_bexp__196 != high_exp__426 | ne_168403 | prod_sign__50);
  assign has_neg_inf__52 = eq_168404 & eq_168405 & x_sign__100 | eq_168406 & eq_168407 & prod_sign__50;
  assign and_reduce_168506 = &result_exp__165[7:0];
  assign wide_exponent__213 = wide_exponent__211[8:0] & {9{~wide_exponent__211[9]}};
  assign has_pos_inf__71 = ~(x_bexp__540 != high_exp__457 | ne_168417 | x_sign__136) | ~(prod_bexp__268 != high_exp__458 | ne_168419 | prod_sign__68);
  assign has_neg_inf__71 = eq_168420 & eq_168421 & x_sign__136 | eq_168422 & eq_168423 & prod_sign__68;
  assign is_result_nan__146 = is_result_nan__147 & ne_168472;
  assign has_inf_arg__76 = is_result_nan__147 & x_fraction__541 == result_fraction__729;
  assign and_reduce_168520 = &result_exp__225[7:0];
  assign is_result_nan__31 = eq_168307 & ne_168304 | eq_168309 & ne_168306 | has_pos_inf__15 & has_neg_inf__15;
  assign is_operand_inf__15 = eq_168307 & eq_168308 | eq_168309 & eq_168310;
  assign and_reduce_168533 = &wide_exponent__47[7:0];
  assign is_result_nan__66 = eq_168325 & ne_168322 | eq_168327 & ne_168324 | has_pos_inf__32 & has_neg_inf__32;
  assign is_operand_inf__32 = eq_168325 & eq_168326 | eq_168327 & eq_168328;
  assign and_reduce_168546 = &wide_exponent__98[7:0];
  assign is_result_nan__105 = eq_168343 & ne_168340 | eq_168345 & ne_168342 | has_pos_inf__51 & has_neg_inf__51;
  assign is_operand_inf__51 = eq_168343 & eq_168344 | eq_168345 & eq_168346;
  assign and_reduce_168560 = &wide_exponent__155[7:0];
  assign high_exp__255 = 8'hff;
  assign is_result_nan__144 = eq_168363 & ne_168360 | eq_168365 & ne_168362 | has_pos_inf__70 & has_neg_inf__70;
  assign is_operand_inf__70 = eq_168363 & eq_168364 | eq_168365 & eq_168366;
  assign and_reduce_168576 = &wide_exponent__212[7:0];
  assign high_exp__328 = 8'hff;
  assign is_result_nan__14 = eq_168374 & ne_168371 | eq_168376 & ne_168373 | has_pos_inf__7 & has_neg_inf__7;
  assign is_operand_inf__7 = eq_168374 & eq_168375 | eq_168376 & eq_168377;
  assign and_reduce_168584 = &wide_exponent__21[7:0];
  assign fraction_shift__378 = 3'h3;
  assign fraction_shift__251 = 3'h4;
  assign high_exp__121 = 8'hff;
  assign is_result_nan__67 = eq_168389 & ne_168386 | eq_168391 & ne_168388 | has_pos_inf__33 & has_neg_inf__33;
  assign is_operand_inf__33 = eq_168389 & eq_168390 | eq_168391 & eq_168392;
  assign and_reduce_168595 = &wide_exponent__99[7:0];
  assign fraction_shift__396 = 3'h3;
  assign fraction_shift__286 = 3'h4;
  assign high_exp__186 = 8'hff;
  assign is_result_nan__106 = eq_168404 & ne_168401 | eq_168406 & ne_168403 | has_pos_inf__52 & has_neg_inf__52;
  assign is_operand_inf__52 = eq_168404 & eq_168405 | eq_168406 & eq_168407;
  assign and_reduce_168606 = &wide_exponent__156[7:0];
  assign fraction_shift__414 = 3'h3;
  assign fraction_shift__321 = 3'h4;
  assign is_subnormal__55 = $signed(exp__227) <= $signed(10'h000);
  assign high_exp__253 = 8'hff;
  assign result_exp__167 = is_result_nan__142 | has_inf_arg__73 | result_exp__165[8] | and_reduce_168506 ? high_exp__255 : result_exp__165[7:0];
  assign is_result_nan__145 = eq_168420 & ne_168417 | eq_168422 & ne_168419 | has_pos_inf__71 & has_neg_inf__71;
  assign is_operand_inf__71 = eq_168420 & eq_168421 | eq_168422 & eq_168423;
  assign and_reduce_168619 = &wide_exponent__213[7:0];
  assign fraction_shift__432 = 3'h3;
  assign fraction_shift__356 = 3'h4;
  assign is_subnormal__75 = $signed(exp__309) <= $signed(10'h000);
  assign high_exp__325 = 8'hff;
  assign result_exp__227 = is_result_nan__146 | has_inf_arg__76 | result_exp__225[8] | and_reduce_168520 ? high_exp__328 : result_exp__225[7:0];
  assign fraction_shift__379 = 3'h3;
  assign fraction_shift__252 = 3'h4;
  assign high_exp__122 = 8'hff;
  assign fraction_shift__48 = rounding_carry__15 ? fraction_shift__251 : fraction_shift__378;
  assign result_sign__448 = 1'h0;
  assign result_exponent__16 = is_result_nan__31 | is_operand_inf__15 | wide_exponent__47[8] | and_reduce_168533 ? high_exp__121 : wide_exponent__47[7:0];
  assign fraction_shift__397 = 3'h3;
  assign fraction_shift__287 = 3'h4;
  assign high_exp__187 = 8'hff;
  assign fraction_shift__98 = rounding_carry__32 ? fraction_shift__286 : fraction_shift__396;
  assign result_sign__545 = 1'h0;
  assign result_exponent__32 = is_result_nan__66 | is_operand_inf__32 | wide_exponent__98[8] | and_reduce_168546 ? high_exp__186 : wide_exponent__98[7:0];
  assign fraction_shift__415 = 3'h3;
  assign fraction_shift__322 = 3'h4;
  assign high_exp__254 = 8'hff;
  assign result_exp__168 = {8{is_result_nan__108}};
  assign fraction_shift__155 = rounding_carry__51 ? fraction_shift__321 : fraction_shift__414;
  assign result_sign__645 = 1'h0;
  assign result_exponent__51 = is_result_nan__105 | is_operand_inf__51 | wide_exponent__155[8] | and_reduce_168560 ? high_exp__253 : wide_exponent__155[7:0];
  assign result_sign__646 = 1'h0;
  assign fraction_shift__433 = 3'h3;
  assign fraction_shift__357 = 3'h4;
  assign high_exp__327 = 8'hff;
  assign result_exp__228 = {8{is_result_nan__147}};
  assign fraction_shift__212 = rounding_carry__70 ? fraction_shift__356 : fraction_shift__432;
  assign result_sign__755 = 1'h0;
  assign result_exponent__70 = is_result_nan__144 | is_operand_inf__70 | wide_exponent__212[8] | and_reduce_168576 ? high_exp__325 : wide_exponent__212[7:0];
  assign result_sign__756 = 1'h0;
  assign fraction_shift__21 = rounding_carry__7 ? fraction_shift__252 : fraction_shift__379;
  assign result_sign__449 = 1'h0;
  assign result_exponent__7 = is_result_nan__14 | is_operand_inf__7 | wide_exponent__21[8] | and_reduce_168584 ? high_exp__122 : wide_exponent__21[7:0];
  assign shrl_168675 = rounded_fraction__15 >> fraction_shift__48;
  assign fraction_shift__99 = rounding_carry__33 ? fraction_shift__287 : fraction_shift__397;
  assign result_sign__546 = 1'h0;
  assign result_exponent__33 = is_result_nan__67 | is_operand_inf__33 | wide_exponent__99[8] | and_reduce_168595 ? high_exp__187 : wide_exponent__99[7:0];
  assign shrl_168682 = rounded_fraction__32 >> fraction_shift__98;
  assign fraction_shift__156 = rounding_carry__52 ? fraction_shift__322 : fraction_shift__415;
  assign result_sign__647 = 1'h0;
  assign result_exponent__52 = is_result_nan__106 | is_operand_inf__52 | wide_exponent__156[8] | and_reduce_168606 ? high_exp__254 : wide_exponent__156[7:0];
  assign result_sign__648 = 1'h0;
  assign shrl_168691 = rounded_fraction__51 >> fraction_shift__155;
  assign fraction_shift__213 = rounding_carry__71 ? fraction_shift__357 : fraction_shift__433;
  assign result_sign__757 = 1'h0;
  assign result_exponent__71 = is_result_nan__145 | is_operand_inf__71 | wide_exponent__213[8] | and_reduce_168619 ? high_exp__327 : wide_exponent__213[7:0];
  assign result_sign__758 = 1'h0;
  assign shrl_168702 = rounded_fraction__70 >> fraction_shift__212;
  assign shrl_168707 = rounded_fraction__7 >> fraction_shift__21;
  assign result_fraction__93 = shrl_168675[22:0];
  assign sum__16 = {result_sign__448, result_exponent__16} + concat_162193;
  assign shrl_168713 = rounded_fraction__33 >> fraction_shift__99;
  assign result_fraction__196 = shrl_168682[22:0];
  assign sum__34 = {result_sign__545, result_exponent__32} + concat_165370;
  assign shrl_168719 = rounded_fraction__52 >> fraction_shift__156;
  assign result_fraction__313 = shrl_168691[22:0];
  assign result_fraction__319 = fraction__499[22:0];
  assign sum__53 = {result_sign__645, result_exponent__51} + {result_sign__646, ~result_exp__167};
  assign shrl_168728 = rounded_fraction__71 >> fraction_shift__213;
  assign result_fraction__430 = shrl_168702[22:0];
  assign result_fraction__436 = fraction__678[22:0];
  assign sum__72 = {result_sign__755, result_exponent__70} + {result_sign__756, ~result_exp__227};
  assign result_fraction__40 = shrl_168707[22:0];
  assign sum__8 = {result_sign__449, result_exponent__7} + concat_162166;
  assign result_fraction__94 = result_fraction__93 & {23{~(is_operand_inf__15 | wide_exponent__47[8] | and_reduce_168533 | ~((|wide_exponent__47[8:1]) | wide_exponent__47[0]))}};
  assign nan_fraction__96 = 23'h40_0000;
  assign result_fraction__197 = shrl_168713[22:0];
  assign sum__35 = {result_sign__546, result_exponent__33} + concat_163691;
  assign result_fraction__198 = result_fraction__196 & {23{~(is_operand_inf__32 | wide_exponent__98[8] | and_reduce_168546 | ~((|wide_exponent__98[8:1]) | wide_exponent__98[0]))}};
  assign nan_fraction__123 = 23'h40_0000;
  assign result_fraction__314 = shrl_168719[22:0];
  assign sum__54 = {result_sign__647, result_exponent__52} + {result_sign__648, ~result_exp__168};
  assign result_fraction__315 = result_fraction__313 & {23{~(is_operand_inf__51 | wide_exponent__155[8] | and_reduce_168560 | ~((|wide_exponent__155[8:1]) | wide_exponent__155[0]))}};
  assign nan_fraction__151 = 23'h40_0000;
  assign result_fraction__321 = result_fraction__319 & {23{~(has_inf_arg__73 | result_exp__165[8] | and_reduce_168506 | is_subnormal__55)}};
  assign nan_fraction__153 = 23'h40_0000;
  assign result_fraction__431 = shrl_168728[22:0];
  assign sum__73 = {result_sign__757, result_exponent__71} + {result_sign__758, ~result_exp__228};
  assign result_fraction__432 = result_fraction__430 & {23{~(is_operand_inf__70 | wide_exponent__212[8] | and_reduce_168576 | ~((|wide_exponent__212[8:1]) | wide_exponent__212[0]))}};
  assign nan_fraction__180 = 23'h40_0000;
  assign result_fraction__438 = result_fraction__436 & {23{~(has_inf_arg__76 | result_exp__225[8] | and_reduce_168520 | is_subnormal__75)}};
  assign nan_fraction__182 = 23'h40_0000;
  assign result_fraction__41 = result_fraction__40 & {23{~(is_operand_inf__7 | wide_exponent__21[8] | and_reduce_168584 | ~((|wide_exponent__21[8:1]) | wide_exponent__21[0]))}};
  assign nan_fraction__97 = 23'h40_0000;
  assign result_fraction__95 = is_result_nan__31 ? nan_fraction__96 : result_fraction__94;
  assign prod_bexp__66 = sum__16[8] ? result_exp__204 : result_exponent__16;
  assign x_bexp__779 = 8'h00;
  assign result_fraction__199 = result_fraction__197 & {23{~(is_operand_inf__33 | wide_exponent__99[8] | and_reduce_168595 | ~((|wide_exponent__99[8:1]) | wide_exponent__99[0]))}};
  assign nan_fraction__124 = 23'h40_0000;
  assign result_fraction__200 = is_result_nan__66 ? nan_fraction__123 : result_fraction__198;
  assign prod_bexp__131 = sum__34[8] ? result_exp__156 : result_exponent__32;
  assign x_bexp__780 = 8'h00;
  assign result_fraction__316 = result_fraction__314 & {23{~(is_operand_inf__52 | wide_exponent__156[8] | and_reduce_168606 | ~((|wide_exponent__156[8:1]) | wide_exponent__156[0]))}};
  assign nan_fraction__152 = 23'h40_0000;
  assign result_fraction__317 = is_result_nan__105 ? nan_fraction__151 : result_fraction__315;
  assign result_fraction__323 = is_result_nan__142 ? nan_fraction__153 : result_fraction__321;
  assign prod_bexp__203 = sum__53[8] ? result_exp__167 : result_exponent__51;
  assign x_bexp__781 = 8'h00;
  assign result_fraction__433 = result_fraction__431 & {23{~(is_operand_inf__71 | wide_exponent__213[8] | and_reduce_168619 | ~((|wide_exponent__213[8:1]) | wide_exponent__213[0]))}};
  assign nan_fraction__181 = 23'h40_0000;
  assign result_fraction__434 = is_result_nan__144 ? nan_fraction__180 : result_fraction__432;
  assign result_fraction__440 = is_result_nan__146 ? nan_fraction__182 : result_fraction__438;
  assign prod_bexp__275 = sum__72[8] ? result_exp__227 : result_exponent__70;
  assign x_bexp__782 = 8'h00;
  assign result_fraction__42 = is_result_nan__14 ? nan_fraction__97 : result_fraction__41;
  assign prod_bexp__30 = sum__8[8] ? result_exp__203 : result_exponent__7;
  assign x_bexp__783 = 8'h00;
  assign fraction_is_zero__15 = add_167640 == 26'h000_0000 & xddend_y__15[2:0] == 3'h0;
  assign prod_fraction__48 = sum__16[8] ? result_fraction__393 : result_fraction__95;
  assign incremented_sum__90 = sum__16[7:0] + 8'h01;
  assign result_fraction__201 = is_result_nan__67 ? nan_fraction__124 : result_fraction__199;
  assign prod_bexp__132 = sum__35[8] ? result_exp__209 : result_exponent__33;
  assign x_bexp__784 = 8'h00;
  assign fraction_is_zero__32 = add_167643 == 26'h000_0000 & xddend_y__31[2:0] == 3'h0;
  assign prod_fraction__97 = sum__34[8] ? result_fraction__300 : result_fraction__200;
  assign incremented_sum__108 = sum__34[7:0] + 8'h01;
  assign result_fraction__318 = is_result_nan__106 ? nan_fraction__152 : result_fraction__316;
  assign result_fraction__479 = {is_result_nan__108, 22'h00_0000};
  assign prod_bexp__204 = sum__54[8] ? result_exp__168 : result_exponent__52;
  assign x_bexp__785 = 8'h00;
  assign fraction_is_zero__51 = add_167646 == 26'h000_0000 & xddend_y__49[2:0] == 3'h0;
  assign prod_fraction__151 = sum__53[8] ? result_fraction__323 : result_fraction__317;
  assign incremented_sum__126 = sum__53[7:0] + 8'h01;
  assign result_fraction__435 = is_result_nan__145 ? nan_fraction__181 : result_fraction__433;
  assign result_fraction__480 = {is_result_nan__147, 22'h00_0000};
  assign prod_bexp__276 = sum__73[8] ? result_exp__228 : result_exponent__71;
  assign x_bexp__786 = 8'h00;
  assign fraction_is_zero__70 = add_167649 == 26'h000_0000 & xddend_y__67[2:0] == 3'h0;
  assign prod_fraction__205 = sum__72[8] ? result_fraction__440 : result_fraction__434;
  assign incremented_sum__144 = sum__72[7:0] + 8'h01;
  assign fraction_is_zero__7 = add_167650 == 26'h000_0000 & xddend_y__7[2:0] == 3'h0;
  assign prod_fraction__22 = sum__8[8] ? result_fraction__475 : result_fraction__42;
  assign incremented_sum__91 = sum__8[7:0] + 8'h01;
  assign wide_y__32 = {2'h1, prod_fraction__48, 3'h0};
  assign x_bexpbs_difference__17 = sum__16[8] ? incremented_sum__90 : ~sum__16[7:0];
  assign fraction_is_zero__33 = add_167653 == 26'h000_0000 & xddend_y__32[2:0] == 3'h0;
  assign prod_fraction__98 = sum__35[8] ? result_fraction__476 : result_fraction__201;
  assign incremented_sum__109 = sum__35[7:0] + 8'h01;
  assign wide_y__67 = {2'h1, prod_fraction__97, 3'h0};
  assign x_bexpbs_difference__33 = sum__34[8] ? incremented_sum__108 : ~sum__34[7:0];
  assign fraction_is_zero__52 = add_167656 == 26'h000_0000 & xddend_y__50[2:0] == 3'h0;
  assign prod_fraction__152 = sum__54[8] ? result_fraction__479 : result_fraction__318;
  assign incremented_sum__127 = sum__54[7:0] + 8'h01;
  assign wide_y__105 = {2'h1, prod_fraction__151, 3'h0};
  assign x_bexpbs_difference__51 = sum__53[8] ? incremented_sum__126 : ~sum__53[7:0];
  assign fraction_is_zero__71 = add_167659 == 26'h000_0000 & xddend_y__68[2:0] == 3'h0;
  assign prod_fraction__206 = sum__73[8] ? result_fraction__480 : result_fraction__435;
  assign incremented_sum__145 = sum__73[7:0] + 8'h01;
  assign wide_y__143 = {2'h1, prod_fraction__205, 3'h0};
  assign x_bexpbs_difference__69 = sum__72[8] ? incremented_sum__144 : ~sum__72[7:0];
  assign wide_y__15 = {2'h1, prod_fraction__22, 3'h0};
  assign x_bexpbs_difference__8 = sum__8[8] ? incremented_sum__91 : ~sum__8[7:0];
  assign concat_168936 = {~(add_167640[25] | fraction_is_zero__15), add_167640[25], fraction_is_zero__15};
  assign x_bexp__134 = sum__16[8] ? result_exponent__16 : result_exp__204;
  assign x_bexp__787 = 8'h00;
  assign wide_y__33 = wide_y__32 & {28{prod_bexp__66 != x_bexp__779}};
  assign sub_168942 = 8'h1c - x_bexpbs_difference__17;
  assign wide_y__68 = {2'h1, prod_fraction__98, 3'h0};
  assign x_bexpbs_difference__34 = sum__35[8] ? incremented_sum__109 : ~sum__35[7:0];
  assign concat_168948 = {~(add_167643[25] | fraction_is_zero__32), add_167643[25], fraction_is_zero__32};
  assign x_bexp__267 = sum__34[8] ? result_exponent__32 : result_exp__156;
  assign x_bexp__788 = 8'h00;
  assign wide_y__69 = wide_y__67 & {28{prod_bexp__131 != x_bexp__780}};
  assign sub_168954 = 8'h1c - x_bexpbs_difference__33;
  assign wide_y__106 = {2'h1, prod_fraction__152, 3'h0};
  assign x_bexpbs_difference__52 = sum__54[8] ? incremented_sum__127 : ~sum__54[7:0];
  assign concat_168960 = {~(add_167646[25] | fraction_is_zero__51), add_167646[25], fraction_is_zero__51};
  assign x_bexp__411 = sum__53[8] ? result_exponent__51 : result_exp__167;
  assign x_bexp__789 = 8'h00;
  assign wide_y__107 = wide_y__105 & {28{prod_bexp__203 != x_bexp__781}};
  assign sub_168966 = 8'h1c - x_bexpbs_difference__51;
  assign wide_y__144 = {2'h1, prod_fraction__206, 3'h0};
  assign x_bexpbs_difference__70 = sum__73[8] ? incremented_sum__145 : ~sum__73[7:0];
  assign concat_168972 = {~(add_167649[25] | fraction_is_zero__70), add_167649[25], fraction_is_zero__70};
  assign x_bexp__555 = sum__72[8] ? result_exponent__70 : result_exp__227;
  assign x_bexp__790 = 8'h00;
  assign wide_y__145 = wide_y__143 & {28{prod_bexp__275 != x_bexp__782}};
  assign sub_168978 = 8'h1c - x_bexpbs_difference__69;
  assign concat_168979 = {~(add_167650[25] | fraction_is_zero__7), add_167650[25], fraction_is_zero__7};
  assign x_bexp__62 = sum__8[8] ? result_exponent__7 : result_exp__203;
  assign x_bexp__791 = 8'h00;
  assign wide_y__16 = wide_y__15 & {28{prod_bexp__30 != x_bexp__783}};
  assign sub_168985 = 8'h1c - x_bexpbs_difference__8;
  assign result_sign__77 = x_sign__32 & prod_sign__15 & concat_168936[0] | ~prod_sign__15 & concat_168936[1] | prod_sign__15 & concat_168936[2];
  assign x_fraction__134 = sum__16[8] ? result_fraction__95 : result_fraction__393;
  assign dropped__16 = sub_168942 >= 8'h1c ? 28'h000_0000 : wide_y__33 << sub_168942;
  assign concat_168993 = {~(add_167653[25] | fraction_is_zero__33), add_167653[25], fraction_is_zero__33};
  assign x_bexp__268 = sum__35[8] ? result_exponent__33 : result_exp__209;
  assign x_bexp__792 = 8'h00;
  assign wide_y__70 = wide_y__68 & {28{prod_bexp__132 != x_bexp__784}};
  assign sub_168999 = 8'h1c - x_bexpbs_difference__34;
  assign result_sign__162 = x_sign__63 & prod_sign__31 & concat_168948[0] | ~prod_sign__31 & concat_168948[1] | prod_sign__31 & concat_168948[2];
  assign x_fraction__267 = sum__34[8] ? result_fraction__200 : result_fraction__300;
  assign dropped__34 = sub_168954 >= 8'h1c ? 28'h000_0000 : wide_y__69 << sub_168954;
  assign concat_169007 = {~(add_167656[25] | fraction_is_zero__52), add_167656[25], fraction_is_zero__52};
  assign x_bexp__412 = sum__54[8] ? result_exponent__52 : result_exp__168;
  assign x_bexp__793 = 8'h00;
  assign wide_y__108 = wide_y__106 & {28{prod_bexp__204 != x_bexp__785}};
  assign sub_169013 = 8'h1c - x_bexpbs_difference__52;
  assign result_sign__259 = x_sign__99 & prod_sign__49 & concat_168960[0] | ~prod_sign__49 & concat_168960[1] | prod_sign__49 & concat_168960[2];
  assign x_fraction__411 = sum__53[8] ? result_fraction__317 : result_fraction__323;
  assign dropped__53 = sub_168966 >= 8'h1c ? 28'h000_0000 : wide_y__107 << sub_168966;
  assign concat_169021 = {~(add_167659[25] | fraction_is_zero__71), add_167659[25], fraction_is_zero__71};
  assign x_bexp__556 = sum__73[8] ? result_exponent__71 : result_exp__228;
  assign x_bexp__794 = 8'h00;
  assign wide_y__146 = wide_y__144 & {28{prod_bexp__276 != x_bexp__786}};
  assign sub_169027 = 8'h1c - x_bexpbs_difference__70;
  assign result_sign__356 = x_sign__135 & prod_sign__67 & concat_168972[0] | ~prod_sign__67 & concat_168972[1] | prod_sign__67 & concat_168972[2];
  assign x_fraction__555 = sum__72[8] ? result_fraction__434 : result_fraction__440;
  assign dropped__72 = sub_168978 >= 8'h1c ? 28'h000_0000 : wide_y__145 << sub_168978;
  assign result_sign__33 = x_sign__14 & prod_sign__7 & concat_168979[0] | ~prod_sign__7 & concat_168979[1] | prod_sign__7 & concat_168979[2];
  assign x_fraction__62 = sum__8[8] ? result_fraction__42 : result_fraction__475;
  assign dropped__8 = sub_168985 >= 8'h1c ? 28'h000_0000 : wide_y__16 << sub_168985;
  assign result_sign__78 = is_operand_inf__15 ? ~has_pos_inf__15 : result_sign__77;
  assign wide_x__32 = {2'h1, x_fraction__134, 3'h0};
  assign result_sign__163 = x_sign__64 & prod_sign__32 & concat_168993[0] | ~prod_sign__32 & concat_168993[1] | prod_sign__32 & concat_168993[2];
  assign x_fraction__268 = sum__35[8] ? result_fraction__201 : result_fraction__476;
  assign dropped__35 = sub_168999 >= 8'h1c ? 28'h000_0000 : wide_y__70 << sub_168999;
  assign result_sign__164 = is_operand_inf__32 ? ~has_pos_inf__32 : result_sign__162;
  assign wide_x__67 = {2'h1, x_fraction__267, 3'h0};
  assign high_exp__485 = 8'hff;
  assign result_sign__260 = x_sign__100 & prod_sign__50 & concat_169007[0] | ~prod_sign__50 & concat_169007[1] | prod_sign__50 & concat_169007[2];
  assign x_fraction__412 = sum__54[8] ? result_fraction__318 : result_fraction__479;
  assign dropped__54 = sub_169013 >= 8'h1c ? 28'h000_0000 : wide_y__108 << sub_169013;
  assign result_sign__261 = is_operand_inf__51 ? ~has_pos_inf__51 : result_sign__259;
  assign wide_x__105 = {2'h1, x_fraction__411, 3'h0};
  assign high_exp__490 = 8'hff;
  assign result_sign__357 = x_sign__136 & prod_sign__68 & concat_169021[0] | ~prod_sign__68 & concat_169021[1] | prod_sign__68 & concat_169021[2];
  assign x_fraction__556 = sum__73[8] ? result_fraction__435 : result_fraction__480;
  assign dropped__73 = sub_169027 >= 8'h1c ? 28'h000_0000 : wide_y__146 << sub_169027;
  assign x_sign__137 = array_index_167783[31:31];
  assign result_sign__358 = is_operand_inf__70 ? ~has_pos_inf__70 : result_sign__356;
  assign wide_x__143 = {2'h1, x_fraction__555, 3'h0};
  assign result_sign__34 = is_operand_inf__7 ? ~has_pos_inf__7 : result_sign__33;
  assign wide_x__15 = {2'h1, x_fraction__62, 3'h0};
  assign result_sign__79 = ~is_result_nan__31 & result_sign__78;
  assign wide_x__33 = wide_x__32 & {28{x_bexp__134 != x_bexp__787}};
  assign result_sign__165 = is_operand_inf__33 ? ~has_pos_inf__33 : result_sign__163;
  assign wide_x__68 = {2'h1, x_fraction__268, 3'h0};
  assign result_sign__166 = ~is_result_nan__66 & result_sign__164;
  assign wide_x__69 = wide_x__67 & {28{x_bexp__267 != x_bexp__788}};
  assign result_sign__262 = is_operand_inf__52 ? ~has_pos_inf__52 : result_sign__260;
  assign wide_x__106 = {2'h1, x_fraction__412, 3'h0};
  assign result_sign__263 = ~is_result_nan__105 & result_sign__261;
  assign wide_x__107 = wide_x__105 & {28{x_bexp__411 != x_bexp__789}};
  assign result_sign__359 = is_operand_inf__71 ? ~has_pos_inf__71 : result_sign__357;
  assign wide_x__144 = {2'h1, x_fraction__556, 3'h0};
  assign result_sign__364 = ~(is_result_nan__147 & ne_168472) & x_sign__137;
  assign result_sign__360 = ~is_result_nan__144 & result_sign__358;
  assign wide_x__145 = wide_x__143 & {28{x_bexp__555 != x_bexp__790}};
  assign result_sign__35 = ~is_result_nan__14 & result_sign__34;
  assign wide_x__16 = wide_x__15 & {28{x_bexp__62 != x_bexp__791}};
  assign x_sign__34 = sum__16[8] ? result_sign__79 : result_sign__160;
  assign prod_sign__16 = sum__16[8] ? result_sign__160 : result_sign__79;
  assign neg_169140 = -wide_x__33;
  assign sticky__50 = {27'h000_0000, dropped__16[27:3] != 25'h000_0000};
  assign result_sign__167 = ~is_result_nan__67 & result_sign__165;
  assign wide_x__70 = wide_x__68 & {28{x_bexp__268 != x_bexp__792}};
  assign x_sign__67 = sum__34[8] ? result_sign__166 : result_sign__248;
  assign prod_sign__33 = sum__34[8] ? result_sign__248 : result_sign__166;
  assign neg_169149 = -wide_x__69;
  assign sticky__106 = {27'h000_0000, dropped__34[27:3] != 25'h000_0000};
  assign result_sign__268 = x_bexp__525 != high_exp__485 & x_sign__134;
  assign result_sign__264 = ~is_result_nan__106 & result_sign__262;
  assign wide_x__108 = wide_x__106 & {28{x_bexp__412 != x_bexp__793}};
  assign x_sign__103 = sum__53[8] ? result_sign__263 : result_sign__354;
  assign prod_sign__51 = sum__53[8] ? result_sign__354 : result_sign__263;
  assign neg_169159 = -wide_x__107;
  assign sticky__165 = {27'h000_0000, dropped__53[27:3] != 25'h000_0000};
  assign result_sign__365 = x_bexp__541 != high_exp__490 & x_sign__137;
  assign result_sign__361 = ~is_result_nan__145 & result_sign__359;
  assign wide_x__146 = wide_x__144 & {28{x_bexp__556 != x_bexp__794}};
  assign x_sign__139 = sum__72[8] ? result_sign__360 : result_sign__364;
  assign prod_sign__69 = sum__72[8] ? result_sign__364 : result_sign__360;
  assign neg_169169 = -wide_x__145;
  assign sticky__224 = {27'h000_0000, dropped__72[27:3] != 25'h000_0000};
  assign x_sign__16 = sum__8[8] ? result_sign__35 : result_sign__324;
  assign prod_sign__8 = sum__8[8] ? result_sign__324 : result_sign__35;
  assign neg_169174 = -wide_x__16;
  assign sticky__24 = {27'h000_0000, dropped__8[27:3] != 25'h000_0000};
  assign xddend_y__16 = (x_bexpbs_difference__17 >= 8'h1c ? 28'h000_0000 : wide_y__33 >> x_bexpbs_difference__17) | sticky__50;
  assign x_sign__68 = sum__35[8] ? result_sign__167 : result_sign__334;
  assign prod_sign__34 = sum__35[8] ? result_sign__334 : result_sign__167;
  assign neg_169183 = -wide_x__70;
  assign sticky__107 = {27'h000_0000, dropped__35[27:3] != 25'h000_0000};
  assign xddend_y__33 = (x_bexpbs_difference__33 >= 8'h1c ? 28'h000_0000 : wide_y__69 >> x_bexpbs_difference__33) | sticky__106;
  assign x_sign__104 = sum__54[8] ? result_sign__264 : result_sign__268;
  assign prod_sign__52 = sum__54[8] ? result_sign__268 : result_sign__264;
  assign neg_169192 = -wide_x__108;
  assign sticky__166 = {27'h000_0000, dropped__54[27:3] != 25'h000_0000};
  assign xddend_y__51 = (x_bexpbs_difference__51 >= 8'h1c ? 28'h000_0000 : wide_y__107 >> x_bexpbs_difference__51) | sticky__165;
  assign x_sign__140 = sum__73[8] ? result_sign__361 : result_sign__365;
  assign prod_sign__70 = sum__73[8] ? result_sign__365 : result_sign__361;
  assign neg_169201 = -wide_x__146;
  assign sticky__225 = {27'h000_0000, dropped__73[27:3] != 25'h000_0000};
  assign xddend_y__69 = (x_bexpbs_difference__69 >= 8'h1c ? 28'h000_0000 : wide_y__145 >> x_bexpbs_difference__69) | sticky__224;
  assign xddend_y__8 = (x_bexpbs_difference__8 >= 8'h1c ? 28'h000_0000 : wide_y__16 >> x_bexpbs_difference__8) | sticky__24;
  assign sel_169212 = x_sign__34 ^ prod_sign__16 ? neg_169140[27:3] : wide_x__33[27:3];
  assign result_sign__1068 = 1'h0;
  assign xddend_y__34 = (x_bexpbs_difference__34 >= 8'h1c ? 28'h000_0000 : wide_y__70 >> x_bexpbs_difference__34) | sticky__107;
  assign sel_169219 = x_sign__67 ^ prod_sign__33 ? neg_169149[27:3] : wide_x__69[27:3];
  assign result_sign__1069 = 1'h0;
  assign xddend_y__52 = (x_bexpbs_difference__52 >= 8'h1c ? 28'h000_0000 : wide_y__108 >> x_bexpbs_difference__52) | sticky__166;
  assign sel_169226 = x_sign__103 ^ prod_sign__51 ? neg_169159[27:3] : wide_x__107[27:3];
  assign result_sign__1070 = 1'h0;
  assign xddend_y__70 = (x_bexpbs_difference__70 >= 8'h1c ? 28'h000_0000 : wide_y__146 >> x_bexpbs_difference__70) | sticky__225;
  assign sel_169233 = x_sign__139 ^ prod_sign__69 ? neg_169169[27:3] : wide_x__145[27:3];
  assign result_sign__1071 = 1'h0;
  assign sel_169236 = x_sign__16 ^ prod_sign__8 ? neg_169174[27:3] : wide_x__16[27:3];
  assign result_sign__1072 = 1'h0;
  assign sel_169241 = x_sign__68 ^ prod_sign__34 ? neg_169183[27:3] : wide_x__70[27:3];
  assign result_sign__1073 = 1'h0;
  assign sel_169246 = x_sign__104 ^ prod_sign__52 ? neg_169192[27:3] : wide_x__108[27:3];
  assign result_sign__1074 = 1'h0;
  assign sel_169251 = x_sign__140 ^ prod_sign__70 ? neg_169201[27:3] : wide_x__146[27:3];
  assign result_sign__1075 = 1'h0;
  assign add_169258 = {{1{sel_169212[24]}}, sel_169212} + {result_sign__1068, xddend_y__16[27:3]};
  assign add_169261 = {{1{sel_169219[24]}}, sel_169219} + {result_sign__1069, xddend_y__33[27:3]};
  assign add_169264 = {{1{sel_169226[24]}}, sel_169226} + {result_sign__1070, xddend_y__51[27:3]};
  assign add_169267 = {{1{sel_169233[24]}}, sel_169233} + {result_sign__1071, xddend_y__69[27:3]};
  assign add_169268 = {{1{sel_169236[24]}}, sel_169236} + {result_sign__1072, xddend_y__8[27:3]};
  assign add_169271 = {{1{sel_169241[24]}}, sel_169241} + {result_sign__1073, xddend_y__34[27:3]};
  assign add_169274 = {{1{sel_169246[24]}}, sel_169246} + {result_sign__1074, xddend_y__52[27:3]};
  assign add_169277 = {{1{sel_169251[24]}}, sel_169251} + {result_sign__1075, xddend_y__70[27:3]};
  assign concat_169282 = {add_169258[24:0], xddend_y__16[2:0]};
  assign concat_169285 = {add_169261[24:0], xddend_y__33[2:0]};
  assign concat_169288 = {add_169264[24:0], xddend_y__51[2:0]};
  assign concat_169291 = {add_169267[24:0], xddend_y__69[2:0]};
  assign concat_169292 = {add_169268[24:0], xddend_y__8[2:0]};
  assign concat_169295 = {add_169271[24:0], xddend_y__34[2:0]};
  assign concat_169298 = {add_169274[24:0], xddend_y__52[2:0]};
  assign concat_169301 = {add_169277[24:0], xddend_y__70[2:0]};
  assign xbs_fraction__16 = add_169258[25] ? -concat_169282 : concat_169282;
  assign xbs_fraction__33 = add_169261[25] ? -concat_169285 : concat_169285;
  assign xbs_fraction__51 = add_169264[25] ? -concat_169288 : concat_169288;
  assign xbs_fraction__69 = add_169267[25] ? -concat_169291 : concat_169291;
  assign xbs_fraction__8 = add_169268[25] ? -concat_169292 : concat_169292;
  assign reverse_169317 = {xbs_fraction__16[0], xbs_fraction__16[1], xbs_fraction__16[2], xbs_fraction__16[3], xbs_fraction__16[4], xbs_fraction__16[5], xbs_fraction__16[6], xbs_fraction__16[7], xbs_fraction__16[8], xbs_fraction__16[9], xbs_fraction__16[10], xbs_fraction__16[11], xbs_fraction__16[12], xbs_fraction__16[13], xbs_fraction__16[14], xbs_fraction__16[15], xbs_fraction__16[16], xbs_fraction__16[17], xbs_fraction__16[18], xbs_fraction__16[19], xbs_fraction__16[20], xbs_fraction__16[21], xbs_fraction__16[22], xbs_fraction__16[23], xbs_fraction__16[24], xbs_fraction__16[25], xbs_fraction__16[26], xbs_fraction__16[27]};
  assign xbs_fraction__34 = add_169271[25] ? -concat_169295 : concat_169295;
  assign reverse_169319 = {xbs_fraction__33[0], xbs_fraction__33[1], xbs_fraction__33[2], xbs_fraction__33[3], xbs_fraction__33[4], xbs_fraction__33[5], xbs_fraction__33[6], xbs_fraction__33[7], xbs_fraction__33[8], xbs_fraction__33[9], xbs_fraction__33[10], xbs_fraction__33[11], xbs_fraction__33[12], xbs_fraction__33[13], xbs_fraction__33[14], xbs_fraction__33[15], xbs_fraction__33[16], xbs_fraction__33[17], xbs_fraction__33[18], xbs_fraction__33[19], xbs_fraction__33[20], xbs_fraction__33[21], xbs_fraction__33[22], xbs_fraction__33[23], xbs_fraction__33[24], xbs_fraction__33[25], xbs_fraction__33[26], xbs_fraction__33[27]};
  assign xbs_fraction__52 = add_169274[25] ? -concat_169298 : concat_169298;
  assign reverse_169321 = {xbs_fraction__51[0], xbs_fraction__51[1], xbs_fraction__51[2], xbs_fraction__51[3], xbs_fraction__51[4], xbs_fraction__51[5], xbs_fraction__51[6], xbs_fraction__51[7], xbs_fraction__51[8], xbs_fraction__51[9], xbs_fraction__51[10], xbs_fraction__51[11], xbs_fraction__51[12], xbs_fraction__51[13], xbs_fraction__51[14], xbs_fraction__51[15], xbs_fraction__51[16], xbs_fraction__51[17], xbs_fraction__51[18], xbs_fraction__51[19], xbs_fraction__51[20], xbs_fraction__51[21], xbs_fraction__51[22], xbs_fraction__51[23], xbs_fraction__51[24], xbs_fraction__51[25], xbs_fraction__51[26], xbs_fraction__51[27]};
  assign xbs_fraction__70 = add_169277[25] ? -concat_169301 : concat_169301;
  assign reverse_169323 = {xbs_fraction__69[0], xbs_fraction__69[1], xbs_fraction__69[2], xbs_fraction__69[3], xbs_fraction__69[4], xbs_fraction__69[5], xbs_fraction__69[6], xbs_fraction__69[7], xbs_fraction__69[8], xbs_fraction__69[9], xbs_fraction__69[10], xbs_fraction__69[11], xbs_fraction__69[12], xbs_fraction__69[13], xbs_fraction__69[14], xbs_fraction__69[15], xbs_fraction__69[16], xbs_fraction__69[17], xbs_fraction__69[18], xbs_fraction__69[19], xbs_fraction__69[20], xbs_fraction__69[21], xbs_fraction__69[22], xbs_fraction__69[23], xbs_fraction__69[24], xbs_fraction__69[25], xbs_fraction__69[26], xbs_fraction__69[27]};
  assign reverse_169324 = {xbs_fraction__8[0], xbs_fraction__8[1], xbs_fraction__8[2], xbs_fraction__8[3], xbs_fraction__8[4], xbs_fraction__8[5], xbs_fraction__8[6], xbs_fraction__8[7], xbs_fraction__8[8], xbs_fraction__8[9], xbs_fraction__8[10], xbs_fraction__8[11], xbs_fraction__8[12], xbs_fraction__8[13], xbs_fraction__8[14], xbs_fraction__8[15], xbs_fraction__8[16], xbs_fraction__8[17], xbs_fraction__8[18], xbs_fraction__8[19], xbs_fraction__8[20], xbs_fraction__8[21], xbs_fraction__8[22], xbs_fraction__8[23], xbs_fraction__8[24], xbs_fraction__8[25], xbs_fraction__8[26], xbs_fraction__8[27]};
  assign one_hot_169325 = {reverse_169317[27:0] == 28'h000_0000, reverse_169317[27] && reverse_169317[26:0] == 27'h000_0000, reverse_169317[26] && reverse_169317[25:0] == 26'h000_0000, reverse_169317[25] && reverse_169317[24:0] == 25'h000_0000, reverse_169317[24] && reverse_169317[23:0] == 24'h00_0000, reverse_169317[23] && reverse_169317[22:0] == 23'h00_0000, reverse_169317[22] && reverse_169317[21:0] == 22'h00_0000, reverse_169317[21] && reverse_169317[20:0] == 21'h00_0000, reverse_169317[20] && reverse_169317[19:0] == 20'h0_0000, reverse_169317[19] && reverse_169317[18:0] == 19'h0_0000, reverse_169317[18] && reverse_169317[17:0] == 18'h0_0000, reverse_169317[17] && reverse_169317[16:0] == 17'h0_0000, reverse_169317[16] && reverse_169317[15:0] == 16'h0000, reverse_169317[15] && reverse_169317[14:0] == 15'h0000, reverse_169317[14] && reverse_169317[13:0] == 14'h0000, reverse_169317[13] && reverse_169317[12:0] == 13'h0000, reverse_169317[12] && reverse_169317[11:0] == 12'h000, reverse_169317[11] && reverse_169317[10:0] == 11'h000, reverse_169317[10] && reverse_169317[9:0] == 10'h000, reverse_169317[9] && reverse_169317[8:0] == 9'h000, reverse_169317[8] && reverse_169317[7:0] == 8'h00, reverse_169317[7] && reverse_169317[6:0] == 7'h00, reverse_169317[6] && reverse_169317[5:0] == 6'h00, reverse_169317[5] && reverse_169317[4:0] == 5'h00, reverse_169317[4] && reverse_169317[3:0] == 4'h0, reverse_169317[3] && reverse_169317[2:0] == 3'h0, reverse_169317[2] && reverse_169317[1:0] == 2'h0, reverse_169317[1] && !reverse_169317[0], reverse_169317[0]};
  assign reverse_169326 = {xbs_fraction__34[0], xbs_fraction__34[1], xbs_fraction__34[2], xbs_fraction__34[3], xbs_fraction__34[4], xbs_fraction__34[5], xbs_fraction__34[6], xbs_fraction__34[7], xbs_fraction__34[8], xbs_fraction__34[9], xbs_fraction__34[10], xbs_fraction__34[11], xbs_fraction__34[12], xbs_fraction__34[13], xbs_fraction__34[14], xbs_fraction__34[15], xbs_fraction__34[16], xbs_fraction__34[17], xbs_fraction__34[18], xbs_fraction__34[19], xbs_fraction__34[20], xbs_fraction__34[21], xbs_fraction__34[22], xbs_fraction__34[23], xbs_fraction__34[24], xbs_fraction__34[25], xbs_fraction__34[26], xbs_fraction__34[27]};
  assign one_hot_169327 = {reverse_169319[27:0] == 28'h000_0000, reverse_169319[27] && reverse_169319[26:0] == 27'h000_0000, reverse_169319[26] && reverse_169319[25:0] == 26'h000_0000, reverse_169319[25] && reverse_169319[24:0] == 25'h000_0000, reverse_169319[24] && reverse_169319[23:0] == 24'h00_0000, reverse_169319[23] && reverse_169319[22:0] == 23'h00_0000, reverse_169319[22] && reverse_169319[21:0] == 22'h00_0000, reverse_169319[21] && reverse_169319[20:0] == 21'h00_0000, reverse_169319[20] && reverse_169319[19:0] == 20'h0_0000, reverse_169319[19] && reverse_169319[18:0] == 19'h0_0000, reverse_169319[18] && reverse_169319[17:0] == 18'h0_0000, reverse_169319[17] && reverse_169319[16:0] == 17'h0_0000, reverse_169319[16] && reverse_169319[15:0] == 16'h0000, reverse_169319[15] && reverse_169319[14:0] == 15'h0000, reverse_169319[14] && reverse_169319[13:0] == 14'h0000, reverse_169319[13] && reverse_169319[12:0] == 13'h0000, reverse_169319[12] && reverse_169319[11:0] == 12'h000, reverse_169319[11] && reverse_169319[10:0] == 11'h000, reverse_169319[10] && reverse_169319[9:0] == 10'h000, reverse_169319[9] && reverse_169319[8:0] == 9'h000, reverse_169319[8] && reverse_169319[7:0] == 8'h00, reverse_169319[7] && reverse_169319[6:0] == 7'h00, reverse_169319[6] && reverse_169319[5:0] == 6'h00, reverse_169319[5] && reverse_169319[4:0] == 5'h00, reverse_169319[4] && reverse_169319[3:0] == 4'h0, reverse_169319[3] && reverse_169319[2:0] == 3'h0, reverse_169319[2] && reverse_169319[1:0] == 2'h0, reverse_169319[1] && !reverse_169319[0], reverse_169319[0]};
  assign reverse_169328 = {xbs_fraction__52[0], xbs_fraction__52[1], xbs_fraction__52[2], xbs_fraction__52[3], xbs_fraction__52[4], xbs_fraction__52[5], xbs_fraction__52[6], xbs_fraction__52[7], xbs_fraction__52[8], xbs_fraction__52[9], xbs_fraction__52[10], xbs_fraction__52[11], xbs_fraction__52[12], xbs_fraction__52[13], xbs_fraction__52[14], xbs_fraction__52[15], xbs_fraction__52[16], xbs_fraction__52[17], xbs_fraction__52[18], xbs_fraction__52[19], xbs_fraction__52[20], xbs_fraction__52[21], xbs_fraction__52[22], xbs_fraction__52[23], xbs_fraction__52[24], xbs_fraction__52[25], xbs_fraction__52[26], xbs_fraction__52[27]};
  assign one_hot_169329 = {reverse_169321[27:0] == 28'h000_0000, reverse_169321[27] && reverse_169321[26:0] == 27'h000_0000, reverse_169321[26] && reverse_169321[25:0] == 26'h000_0000, reverse_169321[25] && reverse_169321[24:0] == 25'h000_0000, reverse_169321[24] && reverse_169321[23:0] == 24'h00_0000, reverse_169321[23] && reverse_169321[22:0] == 23'h00_0000, reverse_169321[22] && reverse_169321[21:0] == 22'h00_0000, reverse_169321[21] && reverse_169321[20:0] == 21'h00_0000, reverse_169321[20] && reverse_169321[19:0] == 20'h0_0000, reverse_169321[19] && reverse_169321[18:0] == 19'h0_0000, reverse_169321[18] && reverse_169321[17:0] == 18'h0_0000, reverse_169321[17] && reverse_169321[16:0] == 17'h0_0000, reverse_169321[16] && reverse_169321[15:0] == 16'h0000, reverse_169321[15] && reverse_169321[14:0] == 15'h0000, reverse_169321[14] && reverse_169321[13:0] == 14'h0000, reverse_169321[13] && reverse_169321[12:0] == 13'h0000, reverse_169321[12] && reverse_169321[11:0] == 12'h000, reverse_169321[11] && reverse_169321[10:0] == 11'h000, reverse_169321[10] && reverse_169321[9:0] == 10'h000, reverse_169321[9] && reverse_169321[8:0] == 9'h000, reverse_169321[8] && reverse_169321[7:0] == 8'h00, reverse_169321[7] && reverse_169321[6:0] == 7'h00, reverse_169321[6] && reverse_169321[5:0] == 6'h00, reverse_169321[5] && reverse_169321[4:0] == 5'h00, reverse_169321[4] && reverse_169321[3:0] == 4'h0, reverse_169321[3] && reverse_169321[2:0] == 3'h0, reverse_169321[2] && reverse_169321[1:0] == 2'h0, reverse_169321[1] && !reverse_169321[0], reverse_169321[0]};
  assign reverse_169330 = {xbs_fraction__70[0], xbs_fraction__70[1], xbs_fraction__70[2], xbs_fraction__70[3], xbs_fraction__70[4], xbs_fraction__70[5], xbs_fraction__70[6], xbs_fraction__70[7], xbs_fraction__70[8], xbs_fraction__70[9], xbs_fraction__70[10], xbs_fraction__70[11], xbs_fraction__70[12], xbs_fraction__70[13], xbs_fraction__70[14], xbs_fraction__70[15], xbs_fraction__70[16], xbs_fraction__70[17], xbs_fraction__70[18], xbs_fraction__70[19], xbs_fraction__70[20], xbs_fraction__70[21], xbs_fraction__70[22], xbs_fraction__70[23], xbs_fraction__70[24], xbs_fraction__70[25], xbs_fraction__70[26], xbs_fraction__70[27]};
  assign one_hot_169331 = {reverse_169323[27:0] == 28'h000_0000, reverse_169323[27] && reverse_169323[26:0] == 27'h000_0000, reverse_169323[26] && reverse_169323[25:0] == 26'h000_0000, reverse_169323[25] && reverse_169323[24:0] == 25'h000_0000, reverse_169323[24] && reverse_169323[23:0] == 24'h00_0000, reverse_169323[23] && reverse_169323[22:0] == 23'h00_0000, reverse_169323[22] && reverse_169323[21:0] == 22'h00_0000, reverse_169323[21] && reverse_169323[20:0] == 21'h00_0000, reverse_169323[20] && reverse_169323[19:0] == 20'h0_0000, reverse_169323[19] && reverse_169323[18:0] == 19'h0_0000, reverse_169323[18] && reverse_169323[17:0] == 18'h0_0000, reverse_169323[17] && reverse_169323[16:0] == 17'h0_0000, reverse_169323[16] && reverse_169323[15:0] == 16'h0000, reverse_169323[15] && reverse_169323[14:0] == 15'h0000, reverse_169323[14] && reverse_169323[13:0] == 14'h0000, reverse_169323[13] && reverse_169323[12:0] == 13'h0000, reverse_169323[12] && reverse_169323[11:0] == 12'h000, reverse_169323[11] && reverse_169323[10:0] == 11'h000, reverse_169323[10] && reverse_169323[9:0] == 10'h000, reverse_169323[9] && reverse_169323[8:0] == 9'h000, reverse_169323[8] && reverse_169323[7:0] == 8'h00, reverse_169323[7] && reverse_169323[6:0] == 7'h00, reverse_169323[6] && reverse_169323[5:0] == 6'h00, reverse_169323[5] && reverse_169323[4:0] == 5'h00, reverse_169323[4] && reverse_169323[3:0] == 4'h0, reverse_169323[3] && reverse_169323[2:0] == 3'h0, reverse_169323[2] && reverse_169323[1:0] == 2'h0, reverse_169323[1] && !reverse_169323[0], reverse_169323[0]};
  assign one_hot_169332 = {reverse_169324[27:0] == 28'h000_0000, reverse_169324[27] && reverse_169324[26:0] == 27'h000_0000, reverse_169324[26] && reverse_169324[25:0] == 26'h000_0000, reverse_169324[25] && reverse_169324[24:0] == 25'h000_0000, reverse_169324[24] && reverse_169324[23:0] == 24'h00_0000, reverse_169324[23] && reverse_169324[22:0] == 23'h00_0000, reverse_169324[22] && reverse_169324[21:0] == 22'h00_0000, reverse_169324[21] && reverse_169324[20:0] == 21'h00_0000, reverse_169324[20] && reverse_169324[19:0] == 20'h0_0000, reverse_169324[19] && reverse_169324[18:0] == 19'h0_0000, reverse_169324[18] && reverse_169324[17:0] == 18'h0_0000, reverse_169324[17] && reverse_169324[16:0] == 17'h0_0000, reverse_169324[16] && reverse_169324[15:0] == 16'h0000, reverse_169324[15] && reverse_169324[14:0] == 15'h0000, reverse_169324[14] && reverse_169324[13:0] == 14'h0000, reverse_169324[13] && reverse_169324[12:0] == 13'h0000, reverse_169324[12] && reverse_169324[11:0] == 12'h000, reverse_169324[11] && reverse_169324[10:0] == 11'h000, reverse_169324[10] && reverse_169324[9:0] == 10'h000, reverse_169324[9] && reverse_169324[8:0] == 9'h000, reverse_169324[8] && reverse_169324[7:0] == 8'h00, reverse_169324[7] && reverse_169324[6:0] == 7'h00, reverse_169324[6] && reverse_169324[5:0] == 6'h00, reverse_169324[5] && reverse_169324[4:0] == 5'h00, reverse_169324[4] && reverse_169324[3:0] == 4'h0, reverse_169324[3] && reverse_169324[2:0] == 3'h0, reverse_169324[2] && reverse_169324[1:0] == 2'h0, reverse_169324[1] && !reverse_169324[0], reverse_169324[0]};
  assign encode_169333 = {one_hot_169325[16] | one_hot_169325[17] | one_hot_169325[18] | one_hot_169325[19] | one_hot_169325[20] | one_hot_169325[21] | one_hot_169325[22] | one_hot_169325[23] | one_hot_169325[24] | one_hot_169325[25] | one_hot_169325[26] | one_hot_169325[27] | one_hot_169325[28], one_hot_169325[8] | one_hot_169325[9] | one_hot_169325[10] | one_hot_169325[11] | one_hot_169325[12] | one_hot_169325[13] | one_hot_169325[14] | one_hot_169325[15] | one_hot_169325[24] | one_hot_169325[25] | one_hot_169325[26] | one_hot_169325[27] | one_hot_169325[28], one_hot_169325[4] | one_hot_169325[5] | one_hot_169325[6] | one_hot_169325[7] | one_hot_169325[12] | one_hot_169325[13] | one_hot_169325[14] | one_hot_169325[15] | one_hot_169325[20] | one_hot_169325[21] | one_hot_169325[22] | one_hot_169325[23] | one_hot_169325[28], one_hot_169325[2] | one_hot_169325[3] | one_hot_169325[6] | one_hot_169325[7] | one_hot_169325[10] | one_hot_169325[11] | one_hot_169325[14] | one_hot_169325[15] | one_hot_169325[18] | one_hot_169325[19] | one_hot_169325[22] | one_hot_169325[23] | one_hot_169325[26] | one_hot_169325[27], one_hot_169325[1] | one_hot_169325[3] | one_hot_169325[5] | one_hot_169325[7] | one_hot_169325[9] | one_hot_169325[11] | one_hot_169325[13] | one_hot_169325[15] | one_hot_169325[17] | one_hot_169325[19] | one_hot_169325[21] | one_hot_169325[23] | one_hot_169325[25] | one_hot_169325[27]};
  assign one_hot_169334 = {reverse_169326[27:0] == 28'h000_0000, reverse_169326[27] && reverse_169326[26:0] == 27'h000_0000, reverse_169326[26] && reverse_169326[25:0] == 26'h000_0000, reverse_169326[25] && reverse_169326[24:0] == 25'h000_0000, reverse_169326[24] && reverse_169326[23:0] == 24'h00_0000, reverse_169326[23] && reverse_169326[22:0] == 23'h00_0000, reverse_169326[22] && reverse_169326[21:0] == 22'h00_0000, reverse_169326[21] && reverse_169326[20:0] == 21'h00_0000, reverse_169326[20] && reverse_169326[19:0] == 20'h0_0000, reverse_169326[19] && reverse_169326[18:0] == 19'h0_0000, reverse_169326[18] && reverse_169326[17:0] == 18'h0_0000, reverse_169326[17] && reverse_169326[16:0] == 17'h0_0000, reverse_169326[16] && reverse_169326[15:0] == 16'h0000, reverse_169326[15] && reverse_169326[14:0] == 15'h0000, reverse_169326[14] && reverse_169326[13:0] == 14'h0000, reverse_169326[13] && reverse_169326[12:0] == 13'h0000, reverse_169326[12] && reverse_169326[11:0] == 12'h000, reverse_169326[11] && reverse_169326[10:0] == 11'h000, reverse_169326[10] && reverse_169326[9:0] == 10'h000, reverse_169326[9] && reverse_169326[8:0] == 9'h000, reverse_169326[8] && reverse_169326[7:0] == 8'h00, reverse_169326[7] && reverse_169326[6:0] == 7'h00, reverse_169326[6] && reverse_169326[5:0] == 6'h00, reverse_169326[5] && reverse_169326[4:0] == 5'h00, reverse_169326[4] && reverse_169326[3:0] == 4'h0, reverse_169326[3] && reverse_169326[2:0] == 3'h0, reverse_169326[2] && reverse_169326[1:0] == 2'h0, reverse_169326[1] && !reverse_169326[0], reverse_169326[0]};
  assign encode_169335 = {one_hot_169327[16] | one_hot_169327[17] | one_hot_169327[18] | one_hot_169327[19] | one_hot_169327[20] | one_hot_169327[21] | one_hot_169327[22] | one_hot_169327[23] | one_hot_169327[24] | one_hot_169327[25] | one_hot_169327[26] | one_hot_169327[27] | one_hot_169327[28], one_hot_169327[8] | one_hot_169327[9] | one_hot_169327[10] | one_hot_169327[11] | one_hot_169327[12] | one_hot_169327[13] | one_hot_169327[14] | one_hot_169327[15] | one_hot_169327[24] | one_hot_169327[25] | one_hot_169327[26] | one_hot_169327[27] | one_hot_169327[28], one_hot_169327[4] | one_hot_169327[5] | one_hot_169327[6] | one_hot_169327[7] | one_hot_169327[12] | one_hot_169327[13] | one_hot_169327[14] | one_hot_169327[15] | one_hot_169327[20] | one_hot_169327[21] | one_hot_169327[22] | one_hot_169327[23] | one_hot_169327[28], one_hot_169327[2] | one_hot_169327[3] | one_hot_169327[6] | one_hot_169327[7] | one_hot_169327[10] | one_hot_169327[11] | one_hot_169327[14] | one_hot_169327[15] | one_hot_169327[18] | one_hot_169327[19] | one_hot_169327[22] | one_hot_169327[23] | one_hot_169327[26] | one_hot_169327[27], one_hot_169327[1] | one_hot_169327[3] | one_hot_169327[5] | one_hot_169327[7] | one_hot_169327[9] | one_hot_169327[11] | one_hot_169327[13] | one_hot_169327[15] | one_hot_169327[17] | one_hot_169327[19] | one_hot_169327[21] | one_hot_169327[23] | one_hot_169327[25] | one_hot_169327[27]};
  assign one_hot_169336 = {reverse_169328[27:0] == 28'h000_0000, reverse_169328[27] && reverse_169328[26:0] == 27'h000_0000, reverse_169328[26] && reverse_169328[25:0] == 26'h000_0000, reverse_169328[25] && reverse_169328[24:0] == 25'h000_0000, reverse_169328[24] && reverse_169328[23:0] == 24'h00_0000, reverse_169328[23] && reverse_169328[22:0] == 23'h00_0000, reverse_169328[22] && reverse_169328[21:0] == 22'h00_0000, reverse_169328[21] && reverse_169328[20:0] == 21'h00_0000, reverse_169328[20] && reverse_169328[19:0] == 20'h0_0000, reverse_169328[19] && reverse_169328[18:0] == 19'h0_0000, reverse_169328[18] && reverse_169328[17:0] == 18'h0_0000, reverse_169328[17] && reverse_169328[16:0] == 17'h0_0000, reverse_169328[16] && reverse_169328[15:0] == 16'h0000, reverse_169328[15] && reverse_169328[14:0] == 15'h0000, reverse_169328[14] && reverse_169328[13:0] == 14'h0000, reverse_169328[13] && reverse_169328[12:0] == 13'h0000, reverse_169328[12] && reverse_169328[11:0] == 12'h000, reverse_169328[11] && reverse_169328[10:0] == 11'h000, reverse_169328[10] && reverse_169328[9:0] == 10'h000, reverse_169328[9] && reverse_169328[8:0] == 9'h000, reverse_169328[8] && reverse_169328[7:0] == 8'h00, reverse_169328[7] && reverse_169328[6:0] == 7'h00, reverse_169328[6] && reverse_169328[5:0] == 6'h00, reverse_169328[5] && reverse_169328[4:0] == 5'h00, reverse_169328[4] && reverse_169328[3:0] == 4'h0, reverse_169328[3] && reverse_169328[2:0] == 3'h0, reverse_169328[2] && reverse_169328[1:0] == 2'h0, reverse_169328[1] && !reverse_169328[0], reverse_169328[0]};
  assign encode_169337 = {one_hot_169329[16] | one_hot_169329[17] | one_hot_169329[18] | one_hot_169329[19] | one_hot_169329[20] | one_hot_169329[21] | one_hot_169329[22] | one_hot_169329[23] | one_hot_169329[24] | one_hot_169329[25] | one_hot_169329[26] | one_hot_169329[27] | one_hot_169329[28], one_hot_169329[8] | one_hot_169329[9] | one_hot_169329[10] | one_hot_169329[11] | one_hot_169329[12] | one_hot_169329[13] | one_hot_169329[14] | one_hot_169329[15] | one_hot_169329[24] | one_hot_169329[25] | one_hot_169329[26] | one_hot_169329[27] | one_hot_169329[28], one_hot_169329[4] | one_hot_169329[5] | one_hot_169329[6] | one_hot_169329[7] | one_hot_169329[12] | one_hot_169329[13] | one_hot_169329[14] | one_hot_169329[15] | one_hot_169329[20] | one_hot_169329[21] | one_hot_169329[22] | one_hot_169329[23] | one_hot_169329[28], one_hot_169329[2] | one_hot_169329[3] | one_hot_169329[6] | one_hot_169329[7] | one_hot_169329[10] | one_hot_169329[11] | one_hot_169329[14] | one_hot_169329[15] | one_hot_169329[18] | one_hot_169329[19] | one_hot_169329[22] | one_hot_169329[23] | one_hot_169329[26] | one_hot_169329[27], one_hot_169329[1] | one_hot_169329[3] | one_hot_169329[5] | one_hot_169329[7] | one_hot_169329[9] | one_hot_169329[11] | one_hot_169329[13] | one_hot_169329[15] | one_hot_169329[17] | one_hot_169329[19] | one_hot_169329[21] | one_hot_169329[23] | one_hot_169329[25] | one_hot_169329[27]};
  assign one_hot_169338 = {reverse_169330[27:0] == 28'h000_0000, reverse_169330[27] && reverse_169330[26:0] == 27'h000_0000, reverse_169330[26] && reverse_169330[25:0] == 26'h000_0000, reverse_169330[25] && reverse_169330[24:0] == 25'h000_0000, reverse_169330[24] && reverse_169330[23:0] == 24'h00_0000, reverse_169330[23] && reverse_169330[22:0] == 23'h00_0000, reverse_169330[22] && reverse_169330[21:0] == 22'h00_0000, reverse_169330[21] && reverse_169330[20:0] == 21'h00_0000, reverse_169330[20] && reverse_169330[19:0] == 20'h0_0000, reverse_169330[19] && reverse_169330[18:0] == 19'h0_0000, reverse_169330[18] && reverse_169330[17:0] == 18'h0_0000, reverse_169330[17] && reverse_169330[16:0] == 17'h0_0000, reverse_169330[16] && reverse_169330[15:0] == 16'h0000, reverse_169330[15] && reverse_169330[14:0] == 15'h0000, reverse_169330[14] && reverse_169330[13:0] == 14'h0000, reverse_169330[13] && reverse_169330[12:0] == 13'h0000, reverse_169330[12] && reverse_169330[11:0] == 12'h000, reverse_169330[11] && reverse_169330[10:0] == 11'h000, reverse_169330[10] && reverse_169330[9:0] == 10'h000, reverse_169330[9] && reverse_169330[8:0] == 9'h000, reverse_169330[8] && reverse_169330[7:0] == 8'h00, reverse_169330[7] && reverse_169330[6:0] == 7'h00, reverse_169330[6] && reverse_169330[5:0] == 6'h00, reverse_169330[5] && reverse_169330[4:0] == 5'h00, reverse_169330[4] && reverse_169330[3:0] == 4'h0, reverse_169330[3] && reverse_169330[2:0] == 3'h0, reverse_169330[2] && reverse_169330[1:0] == 2'h0, reverse_169330[1] && !reverse_169330[0], reverse_169330[0]};
  assign encode_169339 = {one_hot_169331[16] | one_hot_169331[17] | one_hot_169331[18] | one_hot_169331[19] | one_hot_169331[20] | one_hot_169331[21] | one_hot_169331[22] | one_hot_169331[23] | one_hot_169331[24] | one_hot_169331[25] | one_hot_169331[26] | one_hot_169331[27] | one_hot_169331[28], one_hot_169331[8] | one_hot_169331[9] | one_hot_169331[10] | one_hot_169331[11] | one_hot_169331[12] | one_hot_169331[13] | one_hot_169331[14] | one_hot_169331[15] | one_hot_169331[24] | one_hot_169331[25] | one_hot_169331[26] | one_hot_169331[27] | one_hot_169331[28], one_hot_169331[4] | one_hot_169331[5] | one_hot_169331[6] | one_hot_169331[7] | one_hot_169331[12] | one_hot_169331[13] | one_hot_169331[14] | one_hot_169331[15] | one_hot_169331[20] | one_hot_169331[21] | one_hot_169331[22] | one_hot_169331[23] | one_hot_169331[28], one_hot_169331[2] | one_hot_169331[3] | one_hot_169331[6] | one_hot_169331[7] | one_hot_169331[10] | one_hot_169331[11] | one_hot_169331[14] | one_hot_169331[15] | one_hot_169331[18] | one_hot_169331[19] | one_hot_169331[22] | one_hot_169331[23] | one_hot_169331[26] | one_hot_169331[27], one_hot_169331[1] | one_hot_169331[3] | one_hot_169331[5] | one_hot_169331[7] | one_hot_169331[9] | one_hot_169331[11] | one_hot_169331[13] | one_hot_169331[15] | one_hot_169331[17] | one_hot_169331[19] | one_hot_169331[21] | one_hot_169331[23] | one_hot_169331[25] | one_hot_169331[27]};
  assign encode_169340 = {one_hot_169332[16] | one_hot_169332[17] | one_hot_169332[18] | one_hot_169332[19] | one_hot_169332[20] | one_hot_169332[21] | one_hot_169332[22] | one_hot_169332[23] | one_hot_169332[24] | one_hot_169332[25] | one_hot_169332[26] | one_hot_169332[27] | one_hot_169332[28], one_hot_169332[8] | one_hot_169332[9] | one_hot_169332[10] | one_hot_169332[11] | one_hot_169332[12] | one_hot_169332[13] | one_hot_169332[14] | one_hot_169332[15] | one_hot_169332[24] | one_hot_169332[25] | one_hot_169332[26] | one_hot_169332[27] | one_hot_169332[28], one_hot_169332[4] | one_hot_169332[5] | one_hot_169332[6] | one_hot_169332[7] | one_hot_169332[12] | one_hot_169332[13] | one_hot_169332[14] | one_hot_169332[15] | one_hot_169332[20] | one_hot_169332[21] | one_hot_169332[22] | one_hot_169332[23] | one_hot_169332[28], one_hot_169332[2] | one_hot_169332[3] | one_hot_169332[6] | one_hot_169332[7] | one_hot_169332[10] | one_hot_169332[11] | one_hot_169332[14] | one_hot_169332[15] | one_hot_169332[18] | one_hot_169332[19] | one_hot_169332[22] | one_hot_169332[23] | one_hot_169332[26] | one_hot_169332[27], one_hot_169332[1] | one_hot_169332[3] | one_hot_169332[5] | one_hot_169332[7] | one_hot_169332[9] | one_hot_169332[11] | one_hot_169332[13] | one_hot_169332[15] | one_hot_169332[17] | one_hot_169332[19] | one_hot_169332[21] | one_hot_169332[23] | one_hot_169332[25] | one_hot_169332[27]};
  assign encode_169342 = {one_hot_169334[16] | one_hot_169334[17] | one_hot_169334[18] | one_hot_169334[19] | one_hot_169334[20] | one_hot_169334[21] | one_hot_169334[22] | one_hot_169334[23] | one_hot_169334[24] | one_hot_169334[25] | one_hot_169334[26] | one_hot_169334[27] | one_hot_169334[28], one_hot_169334[8] | one_hot_169334[9] | one_hot_169334[10] | one_hot_169334[11] | one_hot_169334[12] | one_hot_169334[13] | one_hot_169334[14] | one_hot_169334[15] | one_hot_169334[24] | one_hot_169334[25] | one_hot_169334[26] | one_hot_169334[27] | one_hot_169334[28], one_hot_169334[4] | one_hot_169334[5] | one_hot_169334[6] | one_hot_169334[7] | one_hot_169334[12] | one_hot_169334[13] | one_hot_169334[14] | one_hot_169334[15] | one_hot_169334[20] | one_hot_169334[21] | one_hot_169334[22] | one_hot_169334[23] | one_hot_169334[28], one_hot_169334[2] | one_hot_169334[3] | one_hot_169334[6] | one_hot_169334[7] | one_hot_169334[10] | one_hot_169334[11] | one_hot_169334[14] | one_hot_169334[15] | one_hot_169334[18] | one_hot_169334[19] | one_hot_169334[22] | one_hot_169334[23] | one_hot_169334[26] | one_hot_169334[27], one_hot_169334[1] | one_hot_169334[3] | one_hot_169334[5] | one_hot_169334[7] | one_hot_169334[9] | one_hot_169334[11] | one_hot_169334[13] | one_hot_169334[15] | one_hot_169334[17] | one_hot_169334[19] | one_hot_169334[21] | one_hot_169334[23] | one_hot_169334[25] | one_hot_169334[27]};
  assign encode_169344 = {one_hot_169336[16] | one_hot_169336[17] | one_hot_169336[18] | one_hot_169336[19] | one_hot_169336[20] | one_hot_169336[21] | one_hot_169336[22] | one_hot_169336[23] | one_hot_169336[24] | one_hot_169336[25] | one_hot_169336[26] | one_hot_169336[27] | one_hot_169336[28], one_hot_169336[8] | one_hot_169336[9] | one_hot_169336[10] | one_hot_169336[11] | one_hot_169336[12] | one_hot_169336[13] | one_hot_169336[14] | one_hot_169336[15] | one_hot_169336[24] | one_hot_169336[25] | one_hot_169336[26] | one_hot_169336[27] | one_hot_169336[28], one_hot_169336[4] | one_hot_169336[5] | one_hot_169336[6] | one_hot_169336[7] | one_hot_169336[12] | one_hot_169336[13] | one_hot_169336[14] | one_hot_169336[15] | one_hot_169336[20] | one_hot_169336[21] | one_hot_169336[22] | one_hot_169336[23] | one_hot_169336[28], one_hot_169336[2] | one_hot_169336[3] | one_hot_169336[6] | one_hot_169336[7] | one_hot_169336[10] | one_hot_169336[11] | one_hot_169336[14] | one_hot_169336[15] | one_hot_169336[18] | one_hot_169336[19] | one_hot_169336[22] | one_hot_169336[23] | one_hot_169336[26] | one_hot_169336[27], one_hot_169336[1] | one_hot_169336[3] | one_hot_169336[5] | one_hot_169336[7] | one_hot_169336[9] | one_hot_169336[11] | one_hot_169336[13] | one_hot_169336[15] | one_hot_169336[17] | one_hot_169336[19] | one_hot_169336[21] | one_hot_169336[23] | one_hot_169336[25] | one_hot_169336[27]};
  assign encode_169346 = {one_hot_169338[16] | one_hot_169338[17] | one_hot_169338[18] | one_hot_169338[19] | one_hot_169338[20] | one_hot_169338[21] | one_hot_169338[22] | one_hot_169338[23] | one_hot_169338[24] | one_hot_169338[25] | one_hot_169338[26] | one_hot_169338[27] | one_hot_169338[28], one_hot_169338[8] | one_hot_169338[9] | one_hot_169338[10] | one_hot_169338[11] | one_hot_169338[12] | one_hot_169338[13] | one_hot_169338[14] | one_hot_169338[15] | one_hot_169338[24] | one_hot_169338[25] | one_hot_169338[26] | one_hot_169338[27] | one_hot_169338[28], one_hot_169338[4] | one_hot_169338[5] | one_hot_169338[6] | one_hot_169338[7] | one_hot_169338[12] | one_hot_169338[13] | one_hot_169338[14] | one_hot_169338[15] | one_hot_169338[20] | one_hot_169338[21] | one_hot_169338[22] | one_hot_169338[23] | one_hot_169338[28], one_hot_169338[2] | one_hot_169338[3] | one_hot_169338[6] | one_hot_169338[7] | one_hot_169338[10] | one_hot_169338[11] | one_hot_169338[14] | one_hot_169338[15] | one_hot_169338[18] | one_hot_169338[19] | one_hot_169338[22] | one_hot_169338[23] | one_hot_169338[26] | one_hot_169338[27], one_hot_169338[1] | one_hot_169338[3] | one_hot_169338[5] | one_hot_169338[7] | one_hot_169338[9] | one_hot_169338[11] | one_hot_169338[13] | one_hot_169338[15] | one_hot_169338[17] | one_hot_169338[19] | one_hot_169338[21] | one_hot_169338[23] | one_hot_169338[25] | one_hot_169338[27]};
  assign cancel__17 = |encode_169333[4:1];
  assign carry_bit__16 = xbs_fraction__16[27];
  assign result_fraction__520 = 23'h00_0000;
  assign cancel__34 = |encode_169335[4:1];
  assign carry_bit__34 = xbs_fraction__33[27];
  assign result_fraction__587 = 23'h00_0000;
  assign cancel__53 = |encode_169337[4:1];
  assign carry_bit__53 = xbs_fraction__51[27];
  assign result_fraction__654 = 23'h00_0000;
  assign cancel__72 = |encode_169339[4:1];
  assign carry_bit__72 = xbs_fraction__69[27];
  assign result_fraction__731 = 23'h00_0000;
  assign cancel__8 = |encode_169340[4:1];
  assign carry_bit__8 = xbs_fraction__8[27];
  assign result_fraction__521 = 23'h00_0000;
  assign leading_zeroes__16 = {result_fraction__520, encode_169333};
  assign cancel__35 = |encode_169342[4:1];
  assign carry_bit__35 = xbs_fraction__34[27];
  assign result_fraction__588 = 23'h00_0000;
  assign leading_zeroes__34 = {result_fraction__587, encode_169335};
  assign cancel__54 = |encode_169344[4:1];
  assign carry_bit__54 = xbs_fraction__52[27];
  assign result_fraction__655 = 23'h00_0000;
  assign leading_zeroes__53 = {result_fraction__654, encode_169337};
  assign cancel__73 = |encode_169346[4:1];
  assign carry_bit__73 = xbs_fraction__70[27];
  assign result_fraction__732 = 23'h00_0000;
  assign leading_zeroes__72 = {result_fraction__731, encode_169339};
  assign leading_zeroes__8 = {result_fraction__521, encode_169340};
  assign carry_fraction__32 = xbs_fraction__16[27:1];
  assign add_169413 = leading_zeroes__16 + 28'hfff_ffff;
  assign leading_zeroes__35 = {result_fraction__588, encode_169342};
  assign carry_fraction__67 = xbs_fraction__33[27:1];
  assign add_169426 = leading_zeroes__34 + 28'hfff_ffff;
  assign leading_zeroes__54 = {result_fraction__655, encode_169344};
  assign carry_fraction__105 = xbs_fraction__51[27:1];
  assign add_169439 = leading_zeroes__53 + 28'hfff_ffff;
  assign leading_zeroes__73 = {result_fraction__732, encode_169346};
  assign carry_fraction__143 = xbs_fraction__69[27:1];
  assign add_169452 = leading_zeroes__72 + 28'hfff_ffff;
  assign array_index_169453 = in_img_unflattened[4'hf];
  assign carry_fraction__15 = xbs_fraction__8[27:1];
  assign add_169460 = leading_zeroes__8 + 28'hfff_ffff;
  assign concat_169461 = {~(carry_bit__16 | cancel__17), ~(carry_bit__16 | ~cancel__17), ~(~carry_bit__16 | cancel__17)};
  assign carry_fraction__33 = carry_fraction__32 | {26'h000_0000, xbs_fraction__16[0]};
  assign cancel_fraction__16 = add_169413 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__16[26:0] << add_169413;
  assign result_sign__617 = 1'h0;
  assign carry_fraction__68 = xbs_fraction__34[27:1];
  assign add_169471 = leading_zeroes__35 + 28'hfff_ffff;
  assign concat_169472 = {~(carry_bit__34 | cancel__34), ~(carry_bit__34 | ~cancel__34), ~(~carry_bit__34 | cancel__34)};
  assign carry_fraction__69 = carry_fraction__67 | {26'h000_0000, xbs_fraction__33[0]};
  assign cancel_fraction__34 = add_169426 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__33[26:0] << add_169426;
  assign result_sign__724 = 1'h0;
  assign carry_fraction__106 = xbs_fraction__52[27:1];
  assign add_169482 = leading_zeroes__54 + 28'hfff_ffff;
  assign concat_169483 = {~(carry_bit__53 | cancel__53), ~(carry_bit__53 | ~cancel__53), ~(~carry_bit__53 | cancel__53)};
  assign carry_fraction__107 = carry_fraction__105 | {26'h000_0000, xbs_fraction__51[0]};
  assign cancel_fraction__53 = add_169439 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__51[26:0] << add_169439;
  assign result_sign__748 = 1'h0;
  assign carry_fraction__144 = xbs_fraction__70[27:1];
  assign add_169493 = leading_zeroes__73 + 28'hfff_ffff;
  assign concat_169494 = {~(carry_bit__72 | cancel__72), ~(carry_bit__72 | ~cancel__72), ~(~carry_bit__72 | cancel__72)};
  assign carry_fraction__145 = carry_fraction__143 | {26'h000_0000, xbs_fraction__69[0]};
  assign cancel_fraction__72 = add_169452 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__69[26:0] << add_169452;
  assign result_sign__760 = 1'h0;
  assign x_bexp__557 = array_index_169453[30:23];
  assign concat_169499 = {~(carry_bit__8 | cancel__8), ~(carry_bit__8 | ~cancel__8), ~(~carry_bit__8 | cancel__8)};
  assign carry_fraction__16 = carry_fraction__15 | {26'h000_0000, xbs_fraction__8[0]};
  assign cancel_fraction__8 = add_169460 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__8[26:0] << add_169460;
  assign shifted_fraction__16 = carry_fraction__33 & {27{concat_169461[0]}} | cancel_fraction__16 & {27{concat_169461[1]}} | xbs_fraction__16[26:0] & {27{concat_169461[2]}};
  assign concat_169505 = {~(carry_bit__35 | cancel__35), ~(carry_bit__35 | ~cancel__35), ~(~carry_bit__35 | cancel__35)};
  assign carry_fraction__70 = carry_fraction__68 | {26'h000_0000, xbs_fraction__34[0]};
  assign cancel_fraction__35 = add_169471 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__34[26:0] << add_169471;
  assign shifted_fraction__34 = carry_fraction__69 & {27{concat_169472[0]}} | cancel_fraction__34 & {27{concat_169472[1]}} | xbs_fraction__33[26:0] & {27{concat_169472[2]}};
  assign concat_169511 = {~(carry_bit__54 | cancel__54), ~(carry_bit__54 | ~cancel__54), ~(~carry_bit__54 | cancel__54)};
  assign carry_fraction__108 = carry_fraction__106 | {26'h000_0000, xbs_fraction__52[0]};
  assign cancel_fraction__54 = add_169482 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__52[26:0] << add_169482;
  assign shifted_fraction__53 = carry_fraction__107 & {27{concat_169483[0]}} | cancel_fraction__53 & {27{concat_169483[1]}} | xbs_fraction__51[26:0] & {27{concat_169483[2]}};
  assign concat_169517 = {~(carry_bit__73 | cancel__73), ~(carry_bit__73 | ~cancel__73), ~(~carry_bit__73 | cancel__73)};
  assign carry_fraction__146 = carry_fraction__144 | {26'h000_0000, xbs_fraction__70[0]};
  assign cancel_fraction__73 = add_169493 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__70[26:0] << add_169493;
  assign shifted_fraction__72 = carry_fraction__145 & {27{concat_169494[0]}} | cancel_fraction__72 & {27{concat_169494[1]}} | xbs_fraction__69[26:0] & {27{concat_169494[2]}};
  assign shifted_fraction__8 = carry_fraction__16 & {27{concat_169499[0]}} | cancel_fraction__8 & {27{concat_169499[1]}} | xbs_fraction__8[26:0] & {27{concat_169499[2]}};
  assign result_sign__1076 = 1'h0;
  assign result_sign__452 = 1'h0;
  assign add_169527 = {result_sign__617, x_bexp__503} + 9'h07f;
  assign shifted_fraction__35 = carry_fraction__70 & {27{concat_169505[0]}} | cancel_fraction__35 & {27{concat_169505[1]}} | xbs_fraction__34[26:0] & {27{concat_169505[2]}};
  assign result_sign__1077 = 1'h0;
  assign result_sign__549 = 1'h0;
  assign add_169532 = {result_sign__724, x_bexp__510} + 9'h07f;
  assign shifted_fraction__54 = carry_fraction__108 & {27{concat_169511[0]}} | cancel_fraction__54 & {27{concat_169511[1]}} | xbs_fraction__52[26:0] & {27{concat_169511[2]}};
  assign result_sign__1078 = 1'h0;
  assign result_sign__651 = 1'h0;
  assign add_169537 = {result_sign__748, x_bexp__541} + 9'h07f;
  assign shifted_fraction__73 = carry_fraction__146 & {27{concat_169517[0]}} | cancel_fraction__73 & {27{concat_169517[1]}} | xbs_fraction__70[26:0] & {27{concat_169517[2]}};
  assign result_sign__1079 = 1'h0;
  assign result_sign__763 = 1'h0;
  assign add_169542 = {result_sign__760, x_bexp__557} + 9'h07f;
  assign x_bexp__795 = 8'h00;
  assign result_sign__759 = 1'h0;
  assign x_fraction__557 = array_index_169453[22:0];
  assign result_sign__1080 = 1'h0;
  assign normal_chunk__16 = shifted_fraction__16[2:0];
  assign fraction_shift__253 = 3'h4;
  assign half_way_chunk__16 = shifted_fraction__16[3:2];
  assign result_sign__1081 = 1'h0;
  assign normal_chunk__34 = shifted_fraction__34[2:0];
  assign fraction_shift__288 = 3'h4;
  assign half_way_chunk__34 = shifted_fraction__34[3:2];
  assign result_sign__1082 = 1'h0;
  assign normal_chunk__53 = shifted_fraction__53[2:0];
  assign fraction_shift__323 = 3'h4;
  assign half_way_chunk__53 = shifted_fraction__53[3:2];
  assign result_sign__1083 = 1'h0;
  assign normal_chunk__72 = shifted_fraction__72[2:0];
  assign fraction_shift__358 = 3'h4;
  assign half_way_chunk__72 = shifted_fraction__72[3:2];
  assign ne_169586 = x_bexp__557 != x_bexp__795;
  assign normal_chunk__8 = shifted_fraction__8[2:0];
  assign fraction_shift__254 = 3'h4;
  assign half_way_chunk__8 = shifted_fraction__8[3:2];
  assign result_sign__450 = 1'h0;
  assign add_169598 = {result_sign__1076, shifted_fraction__16[26:3]} + 25'h000_0001;
  assign exp__68 = {result_sign__452, add_169527} + 10'h381;
  assign normal_chunk__35 = shifted_fraction__35[2:0];
  assign fraction_shift__289 = 3'h4;
  assign half_way_chunk__35 = shifted_fraction__35[3:2];
  assign result_sign__547 = 1'h0;
  assign add_169609 = {result_sign__1077, shifted_fraction__34[26:3]} + 25'h000_0001;
  assign exp__147 = {result_sign__549, add_169532} + 10'h381;
  assign normal_chunk__54 = shifted_fraction__54[2:0];
  assign fraction_shift__324 = 3'h4;
  assign half_way_chunk__54 = shifted_fraction__54[3:2];
  assign result_sign__649 = 1'h0;
  assign add_169620 = {result_sign__1078, shifted_fraction__53[26:3]} + 25'h000_0001;
  assign exp__229 = {result_sign__651, add_169537} + 10'h381;
  assign normal_chunk__73 = shifted_fraction__73[2:0];
  assign fraction_shift__359 = 3'h4;
  assign half_way_chunk__73 = shifted_fraction__73[3:2];
  assign result_sign__761 = 1'h0;
  assign add_169631 = {result_sign__1079, shifted_fraction__72[26:3]} + 25'h000_0001;
  assign exp__311 = {result_sign__763, add_169542} + 10'h381;
  assign x_fraction__559 = {result_sign__759, x_fraction__557} | 24'h80_0000;
  assign result_sign__451 = 1'h0;
  assign add_169639 = {result_sign__1080, shifted_fraction__8[26:3]} + 25'h000_0001;
  assign do_round_up__33 = normal_chunk__16 > fraction_shift__253 | half_way_chunk__16 == 2'h3;
  assign exp__69 = exp__68 & sign_ext_164620;
  assign result_sign__548 = 1'h0;
  assign add_169648 = {result_sign__1081, shifted_fraction__35[26:3]} + 25'h000_0001;
  assign do_round_up__70 = normal_chunk__34 > fraction_shift__288 | half_way_chunk__34 == 2'h3;
  assign exp__149 = exp__147 & sign_ext_164631;
  assign result_sign__650 = 1'h0;
  assign add_169657 = {result_sign__1082, shifted_fraction__54[26:3]} + 25'h000_0001;
  assign do_round_up__109 = normal_chunk__53 > fraction_shift__323 | half_way_chunk__53 == 2'h3;
  assign exp__231 = exp__229 & sign_ext_168003;
  assign result_sign__762 = 1'h0;
  assign add_169666 = {result_sign__1083, shifted_fraction__73[26:3]} + 25'h000_0001;
  assign do_round_up__148 = normal_chunk__72 > fraction_shift__358 | half_way_chunk__72 == 2'h3;
  assign exp__313 = exp__311 & {10{ne_169586}};
  assign x_fraction__561 = x_fraction__559 & {24{ne_169586}};
  assign result_sign__826 = 1'h0;
  assign result_sign__827 = 1'h0;
  assign do_round_up__16 = normal_chunk__8 > fraction_shift__254 | half_way_chunk__8 == 2'h3;
  assign rounded_fraction__16 = do_round_up__33 ? {add_169598, normal_chunk__16} : {result_sign__450, shifted_fraction__16};
  assign do_round_up__71 = normal_chunk__35 > fraction_shift__289 | half_way_chunk__35 == 2'h3;
  assign rounded_fraction__34 = do_round_up__70 ? {add_169609, normal_chunk__34} : {result_sign__547, shifted_fraction__34};
  assign do_round_up__110 = normal_chunk__54 > fraction_shift__324 | half_way_chunk__54 == 2'h3;
  assign rounded_fraction__53 = do_round_up__109 ? {add_169620, normal_chunk__53} : {result_sign__649, shifted_fraction__53};
  assign do_round_up__149 = normal_chunk__73 > fraction_shift__359 | half_way_chunk__73 == 2'h3;
  assign rounded_fraction__72 = do_round_up__148 ? {add_169631, normal_chunk__72} : {result_sign__761, shifted_fraction__72};
  assign rounded_fraction__8 = do_round_up__16 ? {add_169639, normal_chunk__8} : {result_sign__451, shifted_fraction__8};
  assign result_sign__453 = 1'h0;
  assign x_bexp__588 = 8'h00;
  assign rounding_carry__16 = rounded_fraction__16[27];
  assign sel_169701 = $signed(exp__69) <= $signed(10'h000) ? concat_164677 : concat_164676;
  assign rounded_fraction__35 = do_round_up__71 ? {add_169648, normal_chunk__35} : {result_sign__548, shifted_fraction__35};
  assign result_sign__550 = 1'h0;
  assign x_bexp__606 = 8'h00;
  assign rounding_carry__34 = rounded_fraction__34[27];
  assign sel_169706 = $signed(exp__149) <= $signed(10'h000) ? concat_164684 : concat_164683;
  assign rounded_fraction__54 = do_round_up__110 ? {add_169657, normal_chunk__54} : {result_sign__650, shifted_fraction__54};
  assign result_sign__652 = 1'h0;
  assign x_bexp__624 = 8'h00;
  assign rounding_carry__53 = rounded_fraction__53[27];
  assign sel_169711 = $signed(exp__231) <= $signed(10'h000) ? concat_168060 : concat_168059;
  assign rounded_fraction__73 = do_round_up__149 ? {add_169666, normal_chunk__73} : {result_sign__762, shifted_fraction__73};
  assign result_sign__764 = 1'h0;
  assign x_bexp__642 = 8'h00;
  assign rounding_carry__72 = rounded_fraction__72[27];
  assign sel_169716 = $signed(exp__313) <= $signed(10'h000) ? {result_sign__827, x_fraction__561} : {x_fraction__561, result_sign__826};
  assign result_sign__454 = 1'h0;
  assign x_bexp__589 = 8'h00;
  assign rounding_carry__8 = rounded_fraction__8[27];
  assign result_sign__933 = 1'h0;
  assign fraction__158 = sel_169701[23:1];
  assign result_sign__551 = 1'h0;
  assign x_bexp__607 = 8'h00;
  assign rounding_carry__35 = rounded_fraction__35[27];
  assign result_sign__939 = 1'h0;
  assign fraction__334 = sel_169706[23:1];
  assign result_sign__653 = 1'h0;
  assign x_bexp__625 = 8'h00;
  assign rounding_carry__54 = rounded_fraction__54[27];
  assign result_sign__947 = 1'h0;
  assign fraction__513 = sel_169711[23:1];
  assign result_sign__765 = 1'h0;
  assign x_bexp__643 = 8'h00;
  assign rounding_carry__73 = rounded_fraction__73[27];
  assign result_sign__955 = 1'h0;
  assign fraction__692 = sel_169716[23:1];
  assign result_sign__455 = 1'h0;
  assign add_169748 = {result_sign__453, x_bexp__134} + {x_bexp__588, rounding_carry__16};
  assign fraction__159 = {result_sign__933, fraction__158};
  assign result_sign__552 = 1'h0;
  assign add_169758 = {result_sign__550, x_bexp__267} + {x_bexp__606, rounding_carry__34};
  assign fraction__336 = {result_sign__939, fraction__334};
  assign result_sign__654 = 1'h0;
  assign add_169768 = {result_sign__652, x_bexp__411} + {x_bexp__624, rounding_carry__53};
  assign fraction__515 = {result_sign__947, fraction__513};
  assign result_sign__766 = 1'h0;
  assign add_169778 = {result_sign__764, x_bexp__555} + {x_bexp__642, rounding_carry__72};
  assign fraction__694 = {result_sign__955, fraction__692};
  assign result_sign__456 = 1'h0;
  assign add_169786 = {result_sign__454, x_bexp__62} + {x_bexp__589, rounding_carry__8};
  assign do_round_up__34 = sel_169701[0] & sel_169701[1];
  assign add_169795 = fraction__159 + 24'h00_0001;
  assign result_sign__553 = 1'h0;
  assign add_169797 = {result_sign__551, x_bexp__268} + {x_bexp__607, rounding_carry__35};
  assign do_round_up__72 = sel_169706[0] & sel_169706[1];
  assign add_169806 = fraction__336 + 24'h00_0001;
  assign result_sign__655 = 1'h0;
  assign add_169808 = {result_sign__653, x_bexp__412} + {x_bexp__625, rounding_carry__54};
  assign do_round_up__111 = sel_169711[0] & sel_169711[1];
  assign add_169817 = fraction__515 + 24'h00_0001;
  assign result_sign__767 = 1'h0;
  assign add_169819 = {result_sign__765, x_bexp__556} + {x_bexp__643, rounding_carry__73};
  assign do_round_up__150 = sel_169716[0] & sel_169716[1];
  assign add_169828 = fraction__694 + 24'h00_0001;
  assign add_169834 = {result_sign__455, add_169748} + 10'h001;
  assign fraction__160 = do_round_up__34 ? add_169795 : fraction__159;
  assign add_169844 = {result_sign__552, add_169758} + 10'h001;
  assign fraction__338 = do_round_up__72 ? add_169806 : fraction__336;
  assign add_169854 = {result_sign__654, add_169768} + 10'h001;
  assign fraction__517 = do_round_up__111 ? add_169817 : fraction__515;
  assign add_169864 = {result_sign__766, add_169778} + 10'h001;
  assign fraction__696 = do_round_up__150 ? add_169828 : fraction__694;
  assign add_169869 = {result_sign__456, add_169786} + 10'h001;
  assign wide_exponent__48 = add_169834 - {5'h00, encode_169333};
  assign add_169875 = exp__69 + 10'h001;
  assign add_169876 = {result_sign__553, add_169797} + 10'h001;
  assign wide_exponent__100 = add_169844 - {5'h00, encode_169335};
  assign add_169882 = exp__149 + 10'h001;
  assign add_169883 = {result_sign__655, add_169808} + 10'h001;
  assign wide_exponent__157 = add_169854 - {5'h00, encode_169337};
  assign add_169889 = exp__231 + 10'h001;
  assign add_169890 = {result_sign__767, add_169819} + 10'h001;
  assign wide_exponent__214 = add_169864 - {5'h00, encode_169339};
  assign add_169896 = exp__313 + 10'h001;
  assign wide_exponent__22 = add_169869 - {5'h00, encode_169340};
  assign wide_exponent__49 = wide_exponent__48 & {10{add_169258 != 26'h000_0000 | xddend_y__16[2:0] != 3'h0}};
  assign exp__71 = fraction__160[23] ? add_169875 : exp__69;
  assign wide_exponent__101 = add_169876 - {5'h00, encode_169342};
  assign wide_exponent__102 = wide_exponent__100 & {10{add_169261 != 26'h000_0000 | xddend_y__33[2:0] != 3'h0}};
  assign exp__153 = fraction__338[23] ? add_169882 : exp__149;
  assign wide_exponent__158 = add_169883 - {5'h00, encode_169344};
  assign wide_exponent__159 = wide_exponent__157 & {10{add_169264 != 26'h000_0000 | xddend_y__51[2:0] != 3'h0}};
  assign exp__235 = fraction__517[23] ? add_169889 : exp__231;
  assign wide_exponent__215 = add_169890 - {5'h00, encode_169346};
  assign wide_exponent__216 = wide_exponent__214 & {10{add_169267 != 26'h000_0000 | xddend_y__69[2:0] != 3'h0}};
  assign exp__317 = fraction__696[23] ? add_169896 : exp__313;
  assign wide_exponent__23 = wide_exponent__22 & {10{add_169268 != 26'h000_0000 | xddend_y__8[2:0] != 3'h0}};
  assign high_exp__377 = 8'hff;
  assign result_fraction__783 = 23'h00_0000;
  assign high_exp__378 = 8'hff;
  assign result_fraction__784 = 23'h00_0000;
  assign high_exp__123 = 8'hff;
  assign result_fraction__522 = 23'h00_0000;
  assign high_exp__124 = 8'hff;
  assign result_fraction__523 = 23'h00_0000;
  assign wide_exponent__103 = wide_exponent__101 & {10{add_169271 != 26'h000_0000 | xddend_y__34[2:0] != 3'h0}};
  assign high_exp__409 = 8'hff;
  assign result_fraction__816 = 23'h00_0000;
  assign high_exp__410 = 8'hff;
  assign result_fraction__817 = 23'h00_0000;
  assign high_exp__188 = 8'hff;
  assign result_fraction__589 = 23'h00_0000;
  assign high_exp__189 = 8'hff;
  assign result_fraction__590 = 23'h00_0000;
  assign wide_exponent__160 = wide_exponent__158 & {10{add_169274 != 26'h000_0000 | xddend_y__52[2:0] != 3'h0}};
  assign high_exp__441 = 8'hff;
  assign result_fraction__849 = 23'h00_0000;
  assign high_exp__442 = 8'hff;
  assign result_fraction__850 = 23'h00_0000;
  assign high_exp__256 = 8'hff;
  assign result_fraction__656 = 23'h00_0000;
  assign high_exp__257 = 8'hff;
  assign result_fraction__657 = 23'h00_0000;
  assign wide_exponent__217 = wide_exponent__215 & {10{add_169277 != 26'h000_0000 | xddend_y__70[2:0] != 3'h0}};
  assign high_exp__473 = 8'hff;
  assign result_fraction__882 = 23'h00_0000;
  assign high_exp__474 = 8'hff;
  assign result_fraction__883 = 23'h00_0000;
  assign high_exp__329 = 8'hff;
  assign result_fraction__733 = 23'h00_0000;
  assign high_exp__330 = 8'hff;
  assign result_fraction__734 = 23'h00_0000;
  assign high_exp__363 = 8'hff;
  assign result_fraction__768 = 23'h00_0000;
  assign high_exp__364 = 8'hff;
  assign result_fraction__769 = 23'h00_0000;
  assign high_exp__125 = 8'hff;
  assign result_fraction__524 = 23'h00_0000;
  assign high_exp__126 = 8'hff;
  assign result_fraction__525 = 23'h00_0000;
  assign ne_169972 = x_fraction__134 != result_fraction__783;
  assign ne_169974 = prod_fraction__48 != result_fraction__784;
  assign eq_169975 = x_bexp__134 == high_exp__123;
  assign eq_169976 = x_fraction__134 == result_fraction__522;
  assign eq_169977 = prod_bexp__66 == high_exp__124;
  assign eq_169978 = prod_fraction__48 == result_fraction__523;
  assign result_exp__51 = exp__71[8:0];
  assign high_exp__395 = 8'hff;
  assign result_fraction__801 = 23'h00_0000;
  assign high_exp__396 = 8'hff;
  assign result_fraction__802 = 23'h00_0000;
  assign high_exp__190 = 8'hff;
  assign result_fraction__591 = 23'h00_0000;
  assign high_exp__191 = 8'hff;
  assign result_fraction__592 = 23'h00_0000;
  assign ne_169992 = x_fraction__267 != result_fraction__816;
  assign ne_169994 = prod_fraction__97 != result_fraction__817;
  assign eq_169995 = x_bexp__267 == high_exp__188;
  assign eq_169996 = x_fraction__267 == result_fraction__589;
  assign eq_169997 = prod_bexp__131 == high_exp__189;
  assign eq_169998 = prod_fraction__97 == result_fraction__590;
  assign result_exp__109 = exp__153[8:0];
  assign high_exp__427 = 8'hff;
  assign result_fraction__834 = 23'h00_0000;
  assign high_exp__428 = 8'hff;
  assign result_fraction__835 = 23'h00_0000;
  assign high_exp__258 = 8'hff;
  assign result_fraction__658 = 23'h00_0000;
  assign high_exp__259 = 8'hff;
  assign result_fraction__659 = 23'h00_0000;
  assign ne_170012 = x_fraction__411 != result_fraction__849;
  assign ne_170014 = prod_fraction__151 != result_fraction__850;
  assign eq_170015 = x_bexp__411 == high_exp__256;
  assign eq_170016 = x_fraction__411 == result_fraction__656;
  assign eq_170017 = prod_bexp__203 == high_exp__257;
  assign eq_170018 = prod_fraction__151 == result_fraction__657;
  assign result_exp__169 = exp__235[8:0];
  assign high_exp__459 = 8'hff;
  assign result_fraction__867 = 23'h00_0000;
  assign high_exp__460 = 8'hff;
  assign result_fraction__868 = 23'h00_0000;
  assign high_exp__331 = 8'hff;
  assign result_fraction__735 = 23'h00_0000;
  assign high_exp__332 = 8'hff;
  assign result_fraction__736 = 23'h00_0000;
  assign ne_170032 = x_fraction__555 != result_fraction__882;
  assign ne_170034 = prod_fraction__205 != result_fraction__883;
  assign eq_170035 = x_bexp__555 == high_exp__329;
  assign eq_170036 = x_fraction__555 == result_fraction__733;
  assign eq_170037 = prod_bexp__275 == high_exp__330;
  assign eq_170038 = prod_fraction__205 == result_fraction__734;
  assign result_exp__229 = exp__317[8:0];
  assign ne_170043 = x_fraction__62 != result_fraction__768;
  assign ne_170045 = prod_fraction__22 != result_fraction__769;
  assign eq_170046 = x_bexp__62 == high_exp__125;
  assign eq_170047 = x_fraction__62 == result_fraction__524;
  assign eq_170048 = prod_bexp__30 == high_exp__126;
  assign eq_170049 = prod_fraction__22 == result_fraction__525;
  assign result_exp__52 = result_exp__51 & {9{$signed(exp__71) > $signed(10'h000)}};
  assign ne_170059 = x_fraction__268 != result_fraction__801;
  assign ne_170061 = prod_fraction__98 != result_fraction__802;
  assign eq_170062 = x_bexp__268 == high_exp__190;
  assign eq_170063 = x_fraction__268 == result_fraction__591;
  assign eq_170064 = prod_bexp__132 == high_exp__191;
  assign eq_170065 = prod_fraction__98 == result_fraction__592;
  assign result_exp__111 = result_exp__109 & {9{$signed(exp__153) > $signed(10'h000)}};
  assign ne_170075 = x_fraction__412 != result_fraction__834;
  assign ne_170077 = prod_fraction__152 != result_fraction__835;
  assign eq_170078 = x_bexp__412 == high_exp__258;
  assign eq_170079 = x_fraction__412 == result_fraction__658;
  assign eq_170080 = prod_bexp__204 == high_exp__259;
  assign eq_170081 = prod_fraction__152 == result_fraction__659;
  assign result_exp__171 = result_exp__169 & {9{$signed(exp__235) > $signed(10'h000)}};
  assign ne_170091 = x_fraction__556 != result_fraction__867;
  assign ne_170093 = prod_fraction__206 != result_fraction__868;
  assign eq_170094 = x_bexp__556 == high_exp__331;
  assign eq_170095 = x_fraction__556 == result_fraction__735;
  assign eq_170096 = prod_bexp__276 == high_exp__332;
  assign eq_170097 = prod_fraction__206 == result_fraction__736;
  assign high_exp__334 = 8'hff;
  assign result_fraction__738 = 23'h00_0000;
  assign result_fraction__737 = 23'h00_0000;
  assign result_exp__231 = result_exp__229 & {9{$signed(exp__317) > $signed(10'h000)}};
  assign wide_exponent__50 = wide_exponent__49[8:0] & {9{~wide_exponent__49[9]}};
  assign has_pos_inf__16 = ~(x_bexp__134 != high_exp__377 | ne_169972 | x_sign__34) | ~(prod_bexp__66 != high_exp__378 | ne_169974 | prod_sign__16);
  assign has_neg_inf__16 = eq_169975 & eq_169976 & x_sign__34 | eq_169977 & eq_169978 & prod_sign__16;
  assign wide_exponent__104 = wide_exponent__102[8:0] & {9{~wide_exponent__102[9]}};
  assign has_pos_inf__34 = ~(x_bexp__267 != high_exp__409 | ne_169992 | x_sign__67) | ~(prod_bexp__131 != high_exp__410 | ne_169994 | prod_sign__33);
  assign has_neg_inf__34 = eq_169995 & eq_169996 & x_sign__67 | eq_169997 & eq_169998 & prod_sign__33;
  assign wide_exponent__161 = wide_exponent__159[8:0] & {9{~wide_exponent__159[9]}};
  assign has_pos_inf__53 = ~(x_bexp__411 != high_exp__441 | ne_170012 | x_sign__103) | ~(prod_bexp__203 != high_exp__442 | ne_170014 | prod_sign__51);
  assign has_neg_inf__53 = eq_170015 & eq_170016 & x_sign__103 | eq_170017 & eq_170018 & prod_sign__51;
  assign wide_exponent__218 = wide_exponent__216[8:0] & {9{~wide_exponent__216[9]}};
  assign has_pos_inf__72 = ~(x_bexp__555 != high_exp__473 | ne_170032 | x_sign__139) | ~(prod_bexp__275 != high_exp__474 | ne_170034 | prod_sign__69);
  assign has_neg_inf__72 = eq_170035 & eq_170036 & x_sign__139 | eq_170037 & eq_170038 & prod_sign__69;
  assign eq_170147 = x_bexp__557 == high_exp__334;
  assign ne_170148 = x_fraction__557 != result_fraction__738;
  assign wide_exponent__24 = wide_exponent__23[8:0] & {9{~wide_exponent__23[9]}};
  assign has_pos_inf__8 = ~(x_bexp__62 != high_exp__363 | ne_170043 | x_sign__16) | ~(prod_bexp__30 != high_exp__364 | ne_170045 | prod_sign__8);
  assign has_neg_inf__8 = eq_170046 & eq_170047 & x_sign__16 | eq_170048 & eq_170049 & prod_sign__8;
  assign and_reduce_170162 = &result_exp__52[7:0];
  assign wide_exponent__105 = wide_exponent__103[8:0] & {9{~wide_exponent__103[9]}};
  assign has_pos_inf__35 = ~(x_bexp__268 != high_exp__395 | ne_170059 | x_sign__68) | ~(prod_bexp__132 != high_exp__396 | ne_170061 | prod_sign__34);
  assign has_neg_inf__35 = eq_170062 & eq_170063 & x_sign__68 | eq_170064 & eq_170065 & prod_sign__34;
  assign and_reduce_170174 = &result_exp__111[7:0];
  assign wide_exponent__162 = wide_exponent__160[8:0] & {9{~wide_exponent__160[9]}};
  assign has_pos_inf__54 = ~(x_bexp__412 != high_exp__427 | ne_170075 | x_sign__104) | ~(prod_bexp__204 != high_exp__428 | ne_170077 | prod_sign__52);
  assign has_neg_inf__54 = eq_170078 & eq_170079 & x_sign__104 | eq_170080 & eq_170081 & prod_sign__52;
  assign and_reduce_170186 = &result_exp__171[7:0];
  assign wide_exponent__219 = wide_exponent__217[8:0] & {9{~wide_exponent__217[9]}};
  assign has_pos_inf__73 = ~(x_bexp__556 != high_exp__459 | ne_170091 | x_sign__140) | ~(prod_bexp__276 != high_exp__460 | ne_170093 | prod_sign__70);
  assign has_neg_inf__73 = eq_170094 & eq_170095 & x_sign__140 | eq_170096 & eq_170097 & prod_sign__70;
  assign is_result_nan__150 = eq_170147 & ne_170148;
  assign has_inf_arg__77 = eq_170147 & x_fraction__557 == result_fraction__737;
  assign and_reduce_170200 = &result_exp__231[7:0];
  assign is_result_nan__33 = eq_169975 & ne_169972 | eq_169977 & ne_169974 | has_pos_inf__16 & has_neg_inf__16;
  assign is_operand_inf__16 = eq_169975 & eq_169976 | eq_169977 & eq_169978;
  assign and_reduce_170214 = &wide_exponent__50[7:0];
  assign high_exp__129 = 8'hff;
  assign is_result_nan__70 = eq_169995 & ne_169992 | eq_169997 & ne_169994 | has_pos_inf__34 & has_neg_inf__34;
  assign is_operand_inf__34 = eq_169995 & eq_169996 | eq_169997 & eq_169998;
  assign and_reduce_170230 = &wide_exponent__104[7:0];
  assign high_exp__194 = 8'hff;
  assign is_result_nan__109 = eq_170015 & ne_170012 | eq_170017 & ne_170014 | has_pos_inf__53 & has_neg_inf__53;
  assign is_operand_inf__53 = eq_170015 & eq_170016 | eq_170017 & eq_170018;
  assign and_reduce_170246 = &wide_exponent__161[7:0];
  assign high_exp__262 = 8'hff;
  assign is_result_nan__148 = eq_170035 & ne_170032 | eq_170037 & ne_170034 | has_pos_inf__72 & has_neg_inf__72;
  assign is_operand_inf__72 = eq_170035 & eq_170036 | eq_170037 & eq_170038;
  assign and_reduce_170262 = &wide_exponent__218[7:0];
  assign high_exp__336 = 8'hff;
  assign is_result_nan__16 = eq_170046 & ne_170043 | eq_170048 & ne_170045 | has_pos_inf__8 & has_neg_inf__8;
  assign is_operand_inf__8 = eq_170046 & eq_170047 | eq_170048 & eq_170049;
  assign and_reduce_170270 = &wide_exponent__24[7:0];
  assign fraction_shift__380 = 3'h3;
  assign fraction_shift__255 = 3'h4;
  assign is_subnormal__17 = $signed(exp__71) <= $signed(10'h000);
  assign high_exp__127 = 8'hff;
  assign result_exp__53 = is_result_nan__100 | has_inf_arg__69 | result_exp__52[8] | and_reduce_170162 ? high_exp__129 : result_exp__52[7:0];
  assign is_result_nan__71 = eq_170062 & ne_170059 | eq_170064 & ne_170061 | has_pos_inf__35 & has_neg_inf__35;
  assign is_operand_inf__35 = eq_170062 & eq_170063 | eq_170064 & eq_170065;
  assign and_reduce_170283 = &wide_exponent__105[7:0];
  assign fraction_shift__398 = 3'h3;
  assign fraction_shift__290 = 3'h4;
  assign is_subnormal__37 = $signed(exp__153) <= $signed(10'h000);
  assign high_exp__192 = 8'hff;
  assign result_exp__113 = is_result_nan__139 | has_inf_arg__71 | result_exp__111[8] | and_reduce_170174 ? high_exp__194 : result_exp__111[7:0];
  assign is_result_nan__110 = eq_170078 & ne_170075 | eq_170080 & ne_170077 | has_pos_inf__54 & has_neg_inf__54;
  assign is_operand_inf__54 = eq_170078 & eq_170079 | eq_170080 & eq_170081;
  assign and_reduce_170296 = &wide_exponent__162[7:0];
  assign fraction_shift__416 = 3'h3;
  assign fraction_shift__325 = 3'h4;
  assign is_subnormal__57 = $signed(exp__235) <= $signed(10'h000);
  assign high_exp__260 = 8'hff;
  assign result_exp__173 = is_result_nan__146 | has_inf_arg__76 | result_exp__171[8] | and_reduce_170186 ? high_exp__262 : result_exp__171[7:0];
  assign is_result_nan__149 = eq_170094 & ne_170091 | eq_170096 & ne_170093 | has_pos_inf__73 & has_neg_inf__73;
  assign is_operand_inf__73 = eq_170094 & eq_170095 | eq_170096 & eq_170097;
  assign and_reduce_170309 = &wide_exponent__219[7:0];
  assign fraction_shift__434 = 3'h3;
  assign fraction_shift__360 = 3'h4;
  assign is_subnormal__77 = $signed(exp__317) <= $signed(10'h000);
  assign high_exp__333 = 8'hff;
  assign result_exp__233 = is_result_nan__150 | has_inf_arg__77 | result_exp__231[8] | and_reduce_170200 ? high_exp__336 : result_exp__231[7:0];
  assign fraction_shift__381 = 3'h3;
  assign fraction_shift__256 = 3'h4;
  assign high_exp__128 = 8'hff;
  assign fraction_shift__51 = rounding_carry__16 ? fraction_shift__255 : fraction_shift__380;
  assign result_sign__457 = 1'h0;
  assign result_exponent__17 = is_result_nan__33 | is_operand_inf__16 | wide_exponent__50[8] | and_reduce_170214 ? high_exp__127 : wide_exponent__50[7:0];
  assign result_sign__458 = 1'h0;
  assign fraction_shift__399 = 3'h3;
  assign fraction_shift__291 = 3'h4;
  assign high_exp__193 = 8'hff;
  assign fraction_shift__104 = rounding_carry__34 ? fraction_shift__290 : fraction_shift__398;
  assign result_sign__554 = 1'h0;
  assign result_exponent__34 = is_result_nan__70 | is_operand_inf__34 | wide_exponent__104[8] | and_reduce_170230 ? high_exp__192 : wide_exponent__104[7:0];
  assign result_sign__555 = 1'h0;
  assign fraction_shift__417 = 3'h3;
  assign fraction_shift__326 = 3'h4;
  assign high_exp__261 = 8'hff;
  assign fraction_shift__161 = rounding_carry__53 ? fraction_shift__325 : fraction_shift__416;
  assign result_sign__656 = 1'h0;
  assign result_exponent__53 = is_result_nan__109 | is_operand_inf__53 | wide_exponent__161[8] | and_reduce_170246 ? high_exp__260 : wide_exponent__161[7:0];
  assign result_sign__657 = 1'h0;
  assign fraction_shift__435 = 3'h3;
  assign fraction_shift__361 = 3'h4;
  assign high_exp__335 = 8'hff;
  assign fraction_shift__218 = rounding_carry__72 ? fraction_shift__360 : fraction_shift__434;
  assign result_sign__768 = 1'h0;
  assign result_exponent__72 = is_result_nan__148 | is_operand_inf__72 | wide_exponent__218[8] | and_reduce_170262 ? high_exp__333 : wide_exponent__218[7:0];
  assign result_sign__769 = 1'h0;
  assign fraction_shift__24 = rounding_carry__8 ? fraction_shift__256 : fraction_shift__381;
  assign result_sign__459 = 1'h0;
  assign result_exponent__8 = is_result_nan__16 | is_operand_inf__8 | wide_exponent__24[8] | and_reduce_170270 ? high_exp__128 : wide_exponent__24[7:0];
  assign shrl_170369 = rounded_fraction__16 >> fraction_shift__51;
  assign concat_170373 = {result_sign__458, ~result_exp__53};
  assign fraction_shift__105 = rounding_carry__35 ? fraction_shift__291 : fraction_shift__399;
  assign result_sign__556 = 1'h0;
  assign result_exponent__35 = is_result_nan__71 | is_operand_inf__35 | wide_exponent__105[8] | and_reduce_170283 ? high_exp__193 : wide_exponent__105[7:0];
  assign shrl_170378 = rounded_fraction__34 >> fraction_shift__104;
  assign concat_170382 = {result_sign__555, ~result_exp__113};
  assign fraction_shift__162 = rounding_carry__54 ? fraction_shift__326 : fraction_shift__417;
  assign result_sign__658 = 1'h0;
  assign result_exponent__54 = is_result_nan__110 | is_operand_inf__54 | wide_exponent__162[8] | and_reduce_170296 ? high_exp__261 : wide_exponent__162[7:0];
  assign shrl_170387 = rounded_fraction__53 >> fraction_shift__161;
  assign concat_170391 = {result_sign__657, ~result_exp__173};
  assign fraction_shift__219 = rounding_carry__73 ? fraction_shift__361 : fraction_shift__435;
  assign result_sign__770 = 1'h0;
  assign result_exponent__73 = is_result_nan__149 | is_operand_inf__73 | wide_exponent__219[8] | and_reduce_170309 ? high_exp__335 : wide_exponent__219[7:0];
  assign shrl_170396 = rounded_fraction__72 >> fraction_shift__218;
  assign concat_170400 = {result_sign__769, ~result_exp__233};
  assign shrl_170401 = rounded_fraction__8 >> fraction_shift__24;
  assign result_fraction__99 = shrl_170369[22:0];
  assign result_fraction__102 = fraction__160[22:0];
  assign sum__17 = {result_sign__457, result_exponent__17} + concat_170373;
  assign shrl_170409 = rounded_fraction__35 >> fraction_shift__105;
  assign result_fraction__208 = shrl_170378[22:0];
  assign result_fraction__214 = fraction__338[22:0];
  assign sum__36 = {result_sign__554, result_exponent__34} + concat_170382;
  assign shrl_170417 = rounded_fraction__54 >> fraction_shift__162;
  assign result_fraction__325 = shrl_170387[22:0];
  assign result_fraction__331 = fraction__517[22:0];
  assign sum__55 = {result_sign__656, result_exponent__53} + concat_170391;
  assign shrl_170425 = rounded_fraction__73 >> fraction_shift__219;
  assign result_fraction__442 = shrl_170396[22:0];
  assign result_fraction__448 = fraction__696[22:0];
  assign sum__74 = {result_sign__768, result_exponent__72} + concat_170400;
  assign result_fraction__46 = shrl_170401[22:0];
  assign sum__18 = {result_sign__459, result_exponent__8} + concat_170373;
  assign result_fraction__100 = result_fraction__99 & {23{~(is_operand_inf__16 | wide_exponent__50[8] | and_reduce_170214 | ~((|wide_exponent__50[8:1]) | wide_exponent__50[0]))}};
  assign nan_fraction__98 = 23'h40_0000;
  assign result_fraction__103 = result_fraction__102 & {23{~(has_inf_arg__69 | result_exp__52[8] | and_reduce_170162 | is_subnormal__17)}};
  assign nan_fraction__100 = 23'h40_0000;
  assign result_fraction__209 = shrl_170409[22:0];
  assign sum__37 = {result_sign__556, result_exponent__35} + concat_170382;
  assign result_fraction__210 = result_fraction__208 & {23{~(is_operand_inf__34 | wide_exponent__104[8] | and_reduce_170230 | ~((|wide_exponent__104[8:1]) | wide_exponent__104[0]))}};
  assign nan_fraction__125 = 23'h40_0000;
  assign result_fraction__216 = result_fraction__214 & {23{~(has_inf_arg__71 | result_exp__111[8] | and_reduce_170174 | is_subnormal__37)}};
  assign nan_fraction__127 = 23'h40_0000;
  assign result_fraction__326 = shrl_170417[22:0];
  assign sum__56 = {result_sign__658, result_exponent__54} + concat_170391;
  assign result_fraction__327 = result_fraction__325 & {23{~(is_operand_inf__53 | wide_exponent__161[8] | and_reduce_170246 | ~((|wide_exponent__161[8:1]) | wide_exponent__161[0]))}};
  assign nan_fraction__154 = 23'h40_0000;
  assign result_fraction__333 = result_fraction__331 & {23{~(has_inf_arg__76 | result_exp__171[8] | and_reduce_170186 | is_subnormal__57)}};
  assign nan_fraction__156 = 23'h40_0000;
  assign result_fraction__443 = shrl_170425[22:0];
  assign sum__75 = {result_sign__770, result_exponent__73} + concat_170400;
  assign result_fraction__444 = result_fraction__442 & {23{~(is_operand_inf__72 | wide_exponent__218[8] | and_reduce_170262 | ~((|wide_exponent__218[8:1]) | wide_exponent__218[0]))}};
  assign nan_fraction__183 = 23'h40_0000;
  assign result_fraction__450 = result_fraction__448 & {23{~(has_inf_arg__77 | result_exp__231[8] | and_reduce_170200 | is_subnormal__77)}};
  assign nan_fraction__185 = 23'h40_0000;
  assign result_fraction__47 = result_fraction__46 & {23{~(is_operand_inf__8 | wide_exponent__24[8] | and_reduce_170270 | ~((|wide_exponent__24[8:1]) | wide_exponent__24[0]))}};
  assign nan_fraction__99 = 23'h40_0000;
  assign result_fraction__101 = is_result_nan__33 ? nan_fraction__98 : result_fraction__100;
  assign result_fraction__104 = is_result_nan__100 ? nan_fraction__100 : result_fraction__103;
  assign prod_bexp__70 = sum__17[8] ? result_exp__53 : result_exponent__17;
  assign x_bexp__796 = 8'h00;
  assign result_fraction__211 = result_fraction__209 & {23{~(is_operand_inf__35 | wide_exponent__105[8] | and_reduce_170283 | ~((|wide_exponent__105[8:1]) | wide_exponent__105[0]))}};
  assign nan_fraction__126 = 23'h40_0000;
  assign result_fraction__212 = is_result_nan__70 ? nan_fraction__125 : result_fraction__210;
  assign result_fraction__218 = is_result_nan__139 ? nan_fraction__127 : result_fraction__216;
  assign prod_bexp__139 = sum__36[8] ? result_exp__113 : result_exponent__34;
  assign x_bexp__797 = 8'h00;
  assign result_fraction__328 = result_fraction__326 & {23{~(is_operand_inf__54 | wide_exponent__162[8] | and_reduce_170296 | ~((|wide_exponent__162[8:1]) | wide_exponent__162[0]))}};
  assign nan_fraction__155 = 23'h40_0000;
  assign result_fraction__329 = is_result_nan__109 ? nan_fraction__154 : result_fraction__327;
  assign result_fraction__335 = is_result_nan__146 ? nan_fraction__156 : result_fraction__333;
  assign prod_bexp__211 = sum__55[8] ? result_exp__173 : result_exponent__53;
  assign x_bexp__798 = 8'h00;
  assign result_fraction__445 = result_fraction__443 & {23{~(is_operand_inf__73 | wide_exponent__219[8] | and_reduce_170309 | ~((|wide_exponent__219[8:1]) | wide_exponent__219[0]))}};
  assign nan_fraction__184 = 23'h40_0000;
  assign result_fraction__446 = is_result_nan__148 ? nan_fraction__183 : result_fraction__444;
  assign result_fraction__452 = is_result_nan__150 ? nan_fraction__185 : result_fraction__450;
  assign prod_bexp__283 = sum__74[8] ? result_exp__233 : result_exponent__72;
  assign x_bexp__799 = 8'h00;
  assign result_fraction__48 = is_result_nan__16 ? nan_fraction__99 : result_fraction__47;
  assign prod_bexp__34 = sum__18[8] ? result_exp__53 : result_exponent__8;
  assign x_bexp__800 = 8'h00;
  assign fraction_is_zero__16 = add_169258 == 26'h000_0000 & xddend_y__16[2:0] == 3'h0;
  assign prod_fraction__51 = sum__17[8] ? result_fraction__104 : result_fraction__101;
  assign incremented_sum__92 = sum__17[7:0] + 8'h01;
  assign result_fraction__213 = is_result_nan__71 ? nan_fraction__126 : result_fraction__211;
  assign prod_bexp__140 = sum__37[8] ? result_exp__113 : result_exponent__35;
  assign x_bexp__801 = 8'h00;
  assign fraction_is_zero__34 = add_169261 == 26'h000_0000 & xddend_y__33[2:0] == 3'h0;
  assign prod_fraction__103 = sum__36[8] ? result_fraction__218 : result_fraction__212;
  assign incremented_sum__110 = sum__36[7:0] + 8'h01;
  assign result_fraction__330 = is_result_nan__110 ? nan_fraction__155 : result_fraction__328;
  assign prod_bexp__212 = sum__56[8] ? result_exp__173 : result_exponent__54;
  assign x_bexp__802 = 8'h00;
  assign fraction_is_zero__53 = add_169264 == 26'h000_0000 & xddend_y__51[2:0] == 3'h0;
  assign prod_fraction__157 = sum__55[8] ? result_fraction__335 : result_fraction__329;
  assign incremented_sum__128 = sum__55[7:0] + 8'h01;
  assign result_fraction__447 = is_result_nan__149 ? nan_fraction__184 : result_fraction__445;
  assign prod_bexp__284 = sum__75[8] ? result_exp__233 : result_exponent__73;
  assign x_bexp__803 = 8'h00;
  assign fraction_is_zero__72 = add_169267 == 26'h000_0000 & xddend_y__69[2:0] == 3'h0;
  assign prod_fraction__211 = sum__74[8] ? result_fraction__452 : result_fraction__446;
  assign incremented_sum__146 = sum__74[7:0] + 8'h01;
  assign fraction_is_zero__8 = add_169268 == 26'h000_0000 & xddend_y__8[2:0] == 3'h0;
  assign prod_fraction__25 = sum__18[8] ? result_fraction__104 : result_fraction__48;
  assign incremented_sum__93 = sum__18[7:0] + 8'h01;
  assign wide_y__34 = {2'h1, prod_fraction__51, 3'h0};
  assign x_bexpbs_difference__18 = sum__17[8] ? incremented_sum__92 : ~sum__17[7:0];
  assign fraction_is_zero__35 = add_169271 == 26'h000_0000 & xddend_y__34[2:0] == 3'h0;
  assign prod_fraction__104 = sum__37[8] ? result_fraction__218 : result_fraction__213;
  assign incremented_sum__111 = sum__37[7:0] + 8'h01;
  assign wide_y__71 = {2'h1, prod_fraction__103, 3'h0};
  assign x_bexpbs_difference__35 = sum__36[8] ? incremented_sum__110 : ~sum__36[7:0];
  assign fraction_is_zero__54 = add_169274 == 26'h000_0000 & xddend_y__52[2:0] == 3'h0;
  assign prod_fraction__158 = sum__56[8] ? result_fraction__335 : result_fraction__330;
  assign incremented_sum__129 = sum__56[7:0] + 8'h01;
  assign wide_y__109 = {2'h1, prod_fraction__157, 3'h0};
  assign x_bexpbs_difference__53 = sum__55[8] ? incremented_sum__128 : ~sum__55[7:0];
  assign fraction_is_zero__73 = add_169277 == 26'h000_0000 & xddend_y__70[2:0] == 3'h0;
  assign prod_fraction__212 = sum__75[8] ? result_fraction__452 : result_fraction__447;
  assign incremented_sum__147 = sum__75[7:0] + 8'h01;
  assign wide_y__147 = {2'h1, prod_fraction__211, 3'h0};
  assign x_bexpbs_difference__71 = sum__74[8] ? incremented_sum__146 : ~sum__74[7:0];
  assign wide_y__17 = {2'h1, prod_fraction__25, 3'h0};
  assign x_bexpbs_difference__9 = sum__18[8] ? incremented_sum__93 : ~sum__18[7:0];
  assign concat_170634 = {~(add_169258[25] | fraction_is_zero__16), add_169258[25], fraction_is_zero__16};
  assign x_bexp__142 = sum__17[8] ? result_exponent__17 : result_exp__53;
  assign x_bexp__804 = 8'h00;
  assign wide_y__35 = wide_y__34 & {28{prod_bexp__70 != x_bexp__796}};
  assign sub_170640 = 8'h1c - x_bexpbs_difference__18;
  assign wide_y__72 = {2'h1, prod_fraction__104, 3'h0};
  assign x_bexpbs_difference__36 = sum__37[8] ? incremented_sum__111 : ~sum__37[7:0];
  assign concat_170646 = {~(add_169261[25] | fraction_is_zero__34), add_169261[25], fraction_is_zero__34};
  assign x_bexp__283 = sum__36[8] ? result_exponent__34 : result_exp__113;
  assign x_bexp__805 = 8'h00;
  assign wide_y__73 = wide_y__71 & {28{prod_bexp__139 != x_bexp__797}};
  assign sub_170652 = 8'h1c - x_bexpbs_difference__35;
  assign wide_y__110 = {2'h1, prod_fraction__158, 3'h0};
  assign x_bexpbs_difference__54 = sum__56[8] ? incremented_sum__129 : ~sum__56[7:0];
  assign concat_170658 = {~(add_169264[25] | fraction_is_zero__53), add_169264[25], fraction_is_zero__53};
  assign x_bexp__427 = sum__55[8] ? result_exponent__53 : result_exp__173;
  assign x_bexp__806 = 8'h00;
  assign wide_y__111 = wide_y__109 & {28{prod_bexp__211 != x_bexp__798}};
  assign sub_170664 = 8'h1c - x_bexpbs_difference__53;
  assign wide_y__148 = {2'h1, prod_fraction__212, 3'h0};
  assign x_bexpbs_difference__72 = sum__75[8] ? incremented_sum__147 : ~sum__75[7:0];
  assign concat_170670 = {~(add_169267[25] | fraction_is_zero__72), add_169267[25], fraction_is_zero__72};
  assign x_bexp__571 = sum__74[8] ? result_exponent__72 : result_exp__233;
  assign x_bexp__807 = 8'h00;
  assign wide_y__149 = wide_y__147 & {28{prod_bexp__283 != x_bexp__799}};
  assign sub_170676 = 8'h1c - x_bexpbs_difference__71;
  assign concat_170677 = {~(add_169268[25] | fraction_is_zero__8), add_169268[25], fraction_is_zero__8};
  assign x_bexp__70 = sum__18[8] ? result_exponent__8 : result_exp__53;
  assign x_bexp__808 = 8'h00;
  assign wide_y__36 = wide_y__17 & {28{prod_bexp__34 != x_bexp__800}};
  assign sub_170683 = 8'h1c - x_bexpbs_difference__9;
  assign result_sign__82 = x_sign__34 & prod_sign__16 & concat_170634[0] | ~prod_sign__16 & concat_170634[1] | prod_sign__16 & concat_170634[2];
  assign x_fraction__142 = sum__17[8] ? result_fraction__101 : result_fraction__104;
  assign dropped__17 = sub_170640 >= 8'h1c ? 28'h000_0000 : wide_y__35 << sub_170640;
  assign concat_170691 = {~(add_169271[25] | fraction_is_zero__35), add_169271[25], fraction_is_zero__35};
  assign x_bexp__284 = sum__37[8] ? result_exponent__35 : result_exp__113;
  assign x_bexp__809 = 8'h00;
  assign wide_y__74 = wide_y__72 & {28{prod_bexp__140 != x_bexp__801}};
  assign sub_170697 = 8'h1c - x_bexpbs_difference__36;
  assign result_sign__172 = x_sign__67 & prod_sign__33 & concat_170646[0] | ~prod_sign__33 & concat_170646[1] | prod_sign__33 & concat_170646[2];
  assign x_fraction__283 = sum__36[8] ? result_fraction__212 : result_fraction__218;
  assign dropped__36 = sub_170652 >= 8'h1c ? 28'h000_0000 : wide_y__73 << sub_170652;
  assign concat_170705 = {~(add_169274[25] | fraction_is_zero__54), add_169274[25], fraction_is_zero__54};
  assign x_bexp__428 = sum__56[8] ? result_exponent__54 : result_exp__173;
  assign x_bexp__810 = 8'h00;
  assign wide_y__112 = wide_y__110 & {28{prod_bexp__212 != x_bexp__802}};
  assign sub_170711 = 8'h1c - x_bexpbs_difference__54;
  assign result_sign__269 = x_sign__103 & prod_sign__51 & concat_170658[0] | ~prod_sign__51 & concat_170658[1] | prod_sign__51 & concat_170658[2];
  assign x_fraction__427 = sum__55[8] ? result_fraction__329 : result_fraction__335;
  assign dropped__55 = sub_170664 >= 8'h1c ? 28'h000_0000 : wide_y__111 << sub_170664;
  assign concat_170719 = {~(add_169277[25] | fraction_is_zero__73), add_169277[25], fraction_is_zero__73};
  assign x_bexp__572 = sum__75[8] ? result_exponent__73 : result_exp__233;
  assign x_bexp__811 = 8'h00;
  assign wide_y__150 = wide_y__148 & {28{prod_bexp__284 != x_bexp__803}};
  assign sub_170725 = 8'h1c - x_bexpbs_difference__72;
  assign result_sign__366 = x_sign__139 & prod_sign__69 & concat_170670[0] | ~prod_sign__69 & concat_170670[1] | prod_sign__69 & concat_170670[2];
  assign x_fraction__571 = sum__74[8] ? result_fraction__446 : result_fraction__452;
  assign dropped__74 = sub_170676 >= 8'h1c ? 28'h000_0000 : wide_y__149 << sub_170676;
  assign result_sign__38 = x_sign__16 & prod_sign__8 & concat_170677[0] | ~prod_sign__8 & concat_170677[1] | prod_sign__8 & concat_170677[2];
  assign x_fraction__70 = sum__18[8] ? result_fraction__48 : result_fraction__104;
  assign dropped__18 = sub_170683 >= 8'h1c ? 28'h000_0000 : wide_y__36 << sub_170683;
  assign result_sign__83 = is_operand_inf__16 ? ~has_pos_inf__16 : result_sign__82;
  assign wide_x__34 = {2'h1, x_fraction__142, 3'h0};
  assign result_sign__173 = x_sign__68 & prod_sign__34 & concat_170691[0] | ~prod_sign__34 & concat_170691[1] | prod_sign__34 & concat_170691[2];
  assign x_fraction__284 = sum__37[8] ? result_fraction__213 : result_fraction__218;
  assign dropped__37 = sub_170697 >= 8'h1c ? 28'h000_0000 : wide_y__74 << sub_170697;
  assign result_sign__174 = is_operand_inf__34 ? ~has_pos_inf__34 : result_sign__172;
  assign wide_x__71 = {2'h1, x_fraction__283, 3'h0};
  assign result_sign__270 = x_sign__104 & prod_sign__52 & concat_170705[0] | ~prod_sign__52 & concat_170705[1] | prod_sign__52 & concat_170705[2];
  assign x_fraction__428 = sum__56[8] ? result_fraction__330 : result_fraction__335;
  assign dropped__56 = sub_170711 >= 8'h1c ? 28'h000_0000 : wide_y__112 << sub_170711;
  assign result_sign__271 = is_operand_inf__53 ? ~has_pos_inf__53 : result_sign__269;
  assign wide_x__109 = {2'h1, x_fraction__427, 3'h0};
  assign result_sign__367 = x_sign__140 & prod_sign__70 & concat_170719[0] | ~prod_sign__70 & concat_170719[1] | prod_sign__70 & concat_170719[2];
  assign x_fraction__572 = sum__75[8] ? result_fraction__447 : result_fraction__452;
  assign dropped__75 = sub_170725 >= 8'h1c ? 28'h000_0000 : wide_y__150 << sub_170725;
  assign x_sign__141 = array_index_169453[31:31];
  assign result_sign__368 = is_operand_inf__72 ? ~has_pos_inf__72 : result_sign__366;
  assign wide_x__147 = {2'h1, x_fraction__571, 3'h0};
  assign result_sign__39 = is_operand_inf__8 ? ~has_pos_inf__8 : result_sign__38;
  assign wide_x__17 = {2'h1, x_fraction__70, 3'h0};
  assign result_sign__84 = ~is_result_nan__33 & result_sign__83;
  assign wide_x__35 = wide_x__34 & {28{x_bexp__142 != x_bexp__804}};
  assign result_sign__175 = is_operand_inf__35 ? ~has_pos_inf__35 : result_sign__173;
  assign wide_x__72 = {2'h1, x_fraction__284, 3'h0};
  assign result_sign__176 = ~is_result_nan__70 & result_sign__174;
  assign wide_x__73 = wide_x__71 & {28{x_bexp__283 != x_bexp__805}};
  assign result_sign__272 = is_operand_inf__54 ? ~has_pos_inf__54 : result_sign__270;
  assign wide_x__110 = {2'h1, x_fraction__428, 3'h0};
  assign result_sign__273 = ~is_result_nan__109 & result_sign__271;
  assign wide_x__111 = wide_x__109 & {28{x_bexp__427 != x_bexp__806}};
  assign result_sign__369 = is_operand_inf__73 ? ~has_pos_inf__73 : result_sign__367;
  assign wide_x__148 = {2'h1, x_fraction__572, 3'h0};
  assign result_sign__374 = ~(eq_170147 & ne_170148) & x_sign__141;
  assign result_sign__370 = ~is_result_nan__148 & result_sign__368;
  assign wide_x__149 = wide_x__147 & {28{x_bexp__571 != x_bexp__807}};
  assign result_sign__40 = ~is_result_nan__16 & result_sign__39;
  assign wide_x__36 = wide_x__17 & {28{x_bexp__70 != x_bexp__808}};
  assign x_sign__36 = sum__17[8] ? result_sign__84 : result_sign__248;
  assign prod_sign__17 = sum__17[8] ? result_sign__248 : result_sign__84;
  assign neg_170834 = -wide_x__35;
  assign sticky__53 = {27'h000_0000, dropped__17[27:3] != 25'h000_0000};
  assign result_sign__177 = ~is_result_nan__71 & result_sign__175;
  assign wide_x__74 = wide_x__72 & {28{x_bexp__284 != x_bexp__809}};
  assign x_sign__71 = sum__36[8] ? result_sign__176 : result_sign__345;
  assign prod_sign__35 = sum__36[8] ? result_sign__345 : result_sign__176;
  assign neg_170843 = -wide_x__73;
  assign sticky__112 = {27'h000_0000, dropped__36[27:3] != 25'h000_0000};
  assign result_sign__274 = ~is_result_nan__110 & result_sign__272;
  assign wide_x__112 = wide_x__110 & {28{x_bexp__428 != x_bexp__810}};
  assign x_sign__107 = sum__55[8] ? result_sign__273 : result_sign__364;
  assign prod_sign__53 = sum__55[8] ? result_sign__364 : result_sign__273;
  assign neg_170852 = -wide_x__111;
  assign sticky__171 = {27'h000_0000, dropped__55[27:3] != 25'h000_0000};
  assign result_sign__371 = ~is_result_nan__149 & result_sign__369;
  assign wide_x__150 = wide_x__148 & {28{x_bexp__572 != x_bexp__811}};
  assign x_sign__143 = sum__74[8] ? result_sign__370 : result_sign__374;
  assign prod_sign__71 = sum__74[8] ? result_sign__374 : result_sign__370;
  assign neg_170861 = -wide_x__149;
  assign sticky__230 = {27'h000_0000, dropped__74[27:3] != 25'h000_0000};
  assign x_sign__18 = sum__18[8] ? result_sign__40 : result_sign__248;
  assign prod_sign__18 = sum__18[8] ? result_sign__248 : result_sign__40;
  assign neg_170866 = -wide_x__36;
  assign sticky__54 = {27'h000_0000, dropped__18[27:3] != 25'h000_0000};
  assign xddend_y__17 = (x_bexpbs_difference__18 >= 8'h1c ? 28'h000_0000 : wide_y__35 >> x_bexpbs_difference__18) | sticky__53;
  assign x_sign__72 = sum__37[8] ? result_sign__177 : result_sign__345;
  assign prod_sign__36 = sum__37[8] ? result_sign__345 : result_sign__177;
  assign neg_170875 = -wide_x__74;
  assign sticky__113 = {27'h000_0000, dropped__37[27:3] != 25'h000_0000};
  assign xddend_y__35 = (x_bexpbs_difference__35 >= 8'h1c ? 28'h000_0000 : wide_y__73 >> x_bexpbs_difference__35) | sticky__112;
  assign x_sign__108 = sum__56[8] ? result_sign__274 : result_sign__364;
  assign prod_sign__54 = sum__56[8] ? result_sign__364 : result_sign__274;
  assign neg_170884 = -wide_x__112;
  assign sticky__172 = {27'h000_0000, dropped__56[27:3] != 25'h000_0000};
  assign xddend_y__53 = (x_bexpbs_difference__53 >= 8'h1c ? 28'h000_0000 : wide_y__111 >> x_bexpbs_difference__53) | sticky__171;
  assign x_sign__144 = sum__75[8] ? result_sign__371 : result_sign__374;
  assign prod_sign__72 = sum__75[8] ? result_sign__374 : result_sign__371;
  assign neg_170893 = -wide_x__150;
  assign sticky__231 = {27'h000_0000, dropped__75[27:3] != 25'h000_0000};
  assign xddend_y__71 = (x_bexpbs_difference__71 >= 8'h1c ? 28'h000_0000 : wide_y__149 >> x_bexpbs_difference__71) | sticky__230;
  assign xddend_y__18 = (x_bexpbs_difference__9 >= 8'h1c ? 28'h000_0000 : wide_y__36 >> x_bexpbs_difference__9) | sticky__54;
  assign sel_170904 = x_sign__36 ^ prod_sign__17 ? neg_170834[27:3] : wide_x__35[27:3];
  assign result_sign__1084 = 1'h0;
  assign xddend_y__36 = (x_bexpbs_difference__36 >= 8'h1c ? 28'h000_0000 : wide_y__74 >> x_bexpbs_difference__36) | sticky__113;
  assign sel_170911 = x_sign__71 ^ prod_sign__35 ? neg_170843[27:3] : wide_x__73[27:3];
  assign result_sign__1085 = 1'h0;
  assign xddend_y__54 = (x_bexpbs_difference__54 >= 8'h1c ? 28'h000_0000 : wide_y__112 >> x_bexpbs_difference__54) | sticky__172;
  assign sel_170918 = x_sign__107 ^ prod_sign__53 ? neg_170852[27:3] : wide_x__111[27:3];
  assign result_sign__1086 = 1'h0;
  assign xddend_y__72 = (x_bexpbs_difference__72 >= 8'h1c ? 28'h000_0000 : wide_y__150 >> x_bexpbs_difference__72) | sticky__231;
  assign sel_170925 = x_sign__143 ^ prod_sign__71 ? neg_170861[27:3] : wide_x__149[27:3];
  assign result_sign__1087 = 1'h0;
  assign sel_170928 = x_sign__18 ^ prod_sign__18 ? neg_170866[27:3] : wide_x__36[27:3];
  assign result_sign__1088 = 1'h0;
  assign sel_170933 = x_sign__72 ^ prod_sign__36 ? neg_170875[27:3] : wide_x__74[27:3];
  assign result_sign__1089 = 1'h0;
  assign sel_170938 = x_sign__108 ^ prod_sign__54 ? neg_170884[27:3] : wide_x__112[27:3];
  assign result_sign__1090 = 1'h0;
  assign sel_170943 = x_sign__144 ^ prod_sign__72 ? neg_170893[27:3] : wide_x__150[27:3];
  assign result_sign__1091 = 1'h0;
  assign add_170950 = {{1{sel_170904[24]}}, sel_170904} + {result_sign__1084, xddend_y__17[27:3]};
  assign add_170953 = {{1{sel_170911[24]}}, sel_170911} + {result_sign__1085, xddend_y__35[27:3]};
  assign add_170956 = {{1{sel_170918[24]}}, sel_170918} + {result_sign__1086, xddend_y__53[27:3]};
  assign add_170959 = {{1{sel_170925[24]}}, sel_170925} + {result_sign__1087, xddend_y__71[27:3]};
  assign add_170960 = {{1{sel_170928[24]}}, sel_170928} + {result_sign__1088, xddend_y__18[27:3]};
  assign add_170963 = {{1{sel_170933[24]}}, sel_170933} + {result_sign__1089, xddend_y__36[27:3]};
  assign add_170966 = {{1{sel_170938[24]}}, sel_170938} + {result_sign__1090, xddend_y__54[27:3]};
  assign add_170969 = {{1{sel_170943[24]}}, sel_170943} + {result_sign__1091, xddend_y__72[27:3]};
  assign concat_170974 = {add_170950[24:0], xddend_y__17[2:0]};
  assign concat_170977 = {add_170953[24:0], xddend_y__35[2:0]};
  assign concat_170980 = {add_170956[24:0], xddend_y__53[2:0]};
  assign concat_170983 = {add_170959[24:0], xddend_y__71[2:0]};
  assign concat_170984 = {add_170960[24:0], xddend_y__18[2:0]};
  assign concat_170987 = {add_170963[24:0], xddend_y__36[2:0]};
  assign concat_170990 = {add_170966[24:0], xddend_y__54[2:0]};
  assign concat_170993 = {add_170969[24:0], xddend_y__72[2:0]};
  assign xbs_fraction__17 = add_170950[25] ? -concat_170974 : concat_170974;
  assign xbs_fraction__35 = add_170953[25] ? -concat_170977 : concat_170977;
  assign xbs_fraction__53 = add_170956[25] ? -concat_170980 : concat_170980;
  assign xbs_fraction__71 = add_170959[25] ? -concat_170983 : concat_170983;
  assign xbs_fraction__18 = add_170960[25] ? -concat_170984 : concat_170984;
  assign reverse_171009 = {xbs_fraction__17[0], xbs_fraction__17[1], xbs_fraction__17[2], xbs_fraction__17[3], xbs_fraction__17[4], xbs_fraction__17[5], xbs_fraction__17[6], xbs_fraction__17[7], xbs_fraction__17[8], xbs_fraction__17[9], xbs_fraction__17[10], xbs_fraction__17[11], xbs_fraction__17[12], xbs_fraction__17[13], xbs_fraction__17[14], xbs_fraction__17[15], xbs_fraction__17[16], xbs_fraction__17[17], xbs_fraction__17[18], xbs_fraction__17[19], xbs_fraction__17[20], xbs_fraction__17[21], xbs_fraction__17[22], xbs_fraction__17[23], xbs_fraction__17[24], xbs_fraction__17[25], xbs_fraction__17[26], xbs_fraction__17[27]};
  assign xbs_fraction__36 = add_170963[25] ? -concat_170987 : concat_170987;
  assign reverse_171011 = {xbs_fraction__35[0], xbs_fraction__35[1], xbs_fraction__35[2], xbs_fraction__35[3], xbs_fraction__35[4], xbs_fraction__35[5], xbs_fraction__35[6], xbs_fraction__35[7], xbs_fraction__35[8], xbs_fraction__35[9], xbs_fraction__35[10], xbs_fraction__35[11], xbs_fraction__35[12], xbs_fraction__35[13], xbs_fraction__35[14], xbs_fraction__35[15], xbs_fraction__35[16], xbs_fraction__35[17], xbs_fraction__35[18], xbs_fraction__35[19], xbs_fraction__35[20], xbs_fraction__35[21], xbs_fraction__35[22], xbs_fraction__35[23], xbs_fraction__35[24], xbs_fraction__35[25], xbs_fraction__35[26], xbs_fraction__35[27]};
  assign xbs_fraction__54 = add_170966[25] ? -concat_170990 : concat_170990;
  assign reverse_171013 = {xbs_fraction__53[0], xbs_fraction__53[1], xbs_fraction__53[2], xbs_fraction__53[3], xbs_fraction__53[4], xbs_fraction__53[5], xbs_fraction__53[6], xbs_fraction__53[7], xbs_fraction__53[8], xbs_fraction__53[9], xbs_fraction__53[10], xbs_fraction__53[11], xbs_fraction__53[12], xbs_fraction__53[13], xbs_fraction__53[14], xbs_fraction__53[15], xbs_fraction__53[16], xbs_fraction__53[17], xbs_fraction__53[18], xbs_fraction__53[19], xbs_fraction__53[20], xbs_fraction__53[21], xbs_fraction__53[22], xbs_fraction__53[23], xbs_fraction__53[24], xbs_fraction__53[25], xbs_fraction__53[26], xbs_fraction__53[27]};
  assign xbs_fraction__72 = add_170969[25] ? -concat_170993 : concat_170993;
  assign reverse_171015 = {xbs_fraction__71[0], xbs_fraction__71[1], xbs_fraction__71[2], xbs_fraction__71[3], xbs_fraction__71[4], xbs_fraction__71[5], xbs_fraction__71[6], xbs_fraction__71[7], xbs_fraction__71[8], xbs_fraction__71[9], xbs_fraction__71[10], xbs_fraction__71[11], xbs_fraction__71[12], xbs_fraction__71[13], xbs_fraction__71[14], xbs_fraction__71[15], xbs_fraction__71[16], xbs_fraction__71[17], xbs_fraction__71[18], xbs_fraction__71[19], xbs_fraction__71[20], xbs_fraction__71[21], xbs_fraction__71[22], xbs_fraction__71[23], xbs_fraction__71[24], xbs_fraction__71[25], xbs_fraction__71[26], xbs_fraction__71[27]};
  assign reverse_171016 = {xbs_fraction__18[0], xbs_fraction__18[1], xbs_fraction__18[2], xbs_fraction__18[3], xbs_fraction__18[4], xbs_fraction__18[5], xbs_fraction__18[6], xbs_fraction__18[7], xbs_fraction__18[8], xbs_fraction__18[9], xbs_fraction__18[10], xbs_fraction__18[11], xbs_fraction__18[12], xbs_fraction__18[13], xbs_fraction__18[14], xbs_fraction__18[15], xbs_fraction__18[16], xbs_fraction__18[17], xbs_fraction__18[18], xbs_fraction__18[19], xbs_fraction__18[20], xbs_fraction__18[21], xbs_fraction__18[22], xbs_fraction__18[23], xbs_fraction__18[24], xbs_fraction__18[25], xbs_fraction__18[26], xbs_fraction__18[27]};
  assign one_hot_171017 = {reverse_171009[27:0] == 28'h000_0000, reverse_171009[27] && reverse_171009[26:0] == 27'h000_0000, reverse_171009[26] && reverse_171009[25:0] == 26'h000_0000, reverse_171009[25] && reverse_171009[24:0] == 25'h000_0000, reverse_171009[24] && reverse_171009[23:0] == 24'h00_0000, reverse_171009[23] && reverse_171009[22:0] == 23'h00_0000, reverse_171009[22] && reverse_171009[21:0] == 22'h00_0000, reverse_171009[21] && reverse_171009[20:0] == 21'h00_0000, reverse_171009[20] && reverse_171009[19:0] == 20'h0_0000, reverse_171009[19] && reverse_171009[18:0] == 19'h0_0000, reverse_171009[18] && reverse_171009[17:0] == 18'h0_0000, reverse_171009[17] && reverse_171009[16:0] == 17'h0_0000, reverse_171009[16] && reverse_171009[15:0] == 16'h0000, reverse_171009[15] && reverse_171009[14:0] == 15'h0000, reverse_171009[14] && reverse_171009[13:0] == 14'h0000, reverse_171009[13] && reverse_171009[12:0] == 13'h0000, reverse_171009[12] && reverse_171009[11:0] == 12'h000, reverse_171009[11] && reverse_171009[10:0] == 11'h000, reverse_171009[10] && reverse_171009[9:0] == 10'h000, reverse_171009[9] && reverse_171009[8:0] == 9'h000, reverse_171009[8] && reverse_171009[7:0] == 8'h00, reverse_171009[7] && reverse_171009[6:0] == 7'h00, reverse_171009[6] && reverse_171009[5:0] == 6'h00, reverse_171009[5] && reverse_171009[4:0] == 5'h00, reverse_171009[4] && reverse_171009[3:0] == 4'h0, reverse_171009[3] && reverse_171009[2:0] == 3'h0, reverse_171009[2] && reverse_171009[1:0] == 2'h0, reverse_171009[1] && !reverse_171009[0], reverse_171009[0]};
  assign reverse_171018 = {xbs_fraction__36[0], xbs_fraction__36[1], xbs_fraction__36[2], xbs_fraction__36[3], xbs_fraction__36[4], xbs_fraction__36[5], xbs_fraction__36[6], xbs_fraction__36[7], xbs_fraction__36[8], xbs_fraction__36[9], xbs_fraction__36[10], xbs_fraction__36[11], xbs_fraction__36[12], xbs_fraction__36[13], xbs_fraction__36[14], xbs_fraction__36[15], xbs_fraction__36[16], xbs_fraction__36[17], xbs_fraction__36[18], xbs_fraction__36[19], xbs_fraction__36[20], xbs_fraction__36[21], xbs_fraction__36[22], xbs_fraction__36[23], xbs_fraction__36[24], xbs_fraction__36[25], xbs_fraction__36[26], xbs_fraction__36[27]};
  assign one_hot_171019 = {reverse_171011[27:0] == 28'h000_0000, reverse_171011[27] && reverse_171011[26:0] == 27'h000_0000, reverse_171011[26] && reverse_171011[25:0] == 26'h000_0000, reverse_171011[25] && reverse_171011[24:0] == 25'h000_0000, reverse_171011[24] && reverse_171011[23:0] == 24'h00_0000, reverse_171011[23] && reverse_171011[22:0] == 23'h00_0000, reverse_171011[22] && reverse_171011[21:0] == 22'h00_0000, reverse_171011[21] && reverse_171011[20:0] == 21'h00_0000, reverse_171011[20] && reverse_171011[19:0] == 20'h0_0000, reverse_171011[19] && reverse_171011[18:0] == 19'h0_0000, reverse_171011[18] && reverse_171011[17:0] == 18'h0_0000, reverse_171011[17] && reverse_171011[16:0] == 17'h0_0000, reverse_171011[16] && reverse_171011[15:0] == 16'h0000, reverse_171011[15] && reverse_171011[14:0] == 15'h0000, reverse_171011[14] && reverse_171011[13:0] == 14'h0000, reverse_171011[13] && reverse_171011[12:0] == 13'h0000, reverse_171011[12] && reverse_171011[11:0] == 12'h000, reverse_171011[11] && reverse_171011[10:0] == 11'h000, reverse_171011[10] && reverse_171011[9:0] == 10'h000, reverse_171011[9] && reverse_171011[8:0] == 9'h000, reverse_171011[8] && reverse_171011[7:0] == 8'h00, reverse_171011[7] && reverse_171011[6:0] == 7'h00, reverse_171011[6] && reverse_171011[5:0] == 6'h00, reverse_171011[5] && reverse_171011[4:0] == 5'h00, reverse_171011[4] && reverse_171011[3:0] == 4'h0, reverse_171011[3] && reverse_171011[2:0] == 3'h0, reverse_171011[2] && reverse_171011[1:0] == 2'h0, reverse_171011[1] && !reverse_171011[0], reverse_171011[0]};
  assign reverse_171020 = {xbs_fraction__54[0], xbs_fraction__54[1], xbs_fraction__54[2], xbs_fraction__54[3], xbs_fraction__54[4], xbs_fraction__54[5], xbs_fraction__54[6], xbs_fraction__54[7], xbs_fraction__54[8], xbs_fraction__54[9], xbs_fraction__54[10], xbs_fraction__54[11], xbs_fraction__54[12], xbs_fraction__54[13], xbs_fraction__54[14], xbs_fraction__54[15], xbs_fraction__54[16], xbs_fraction__54[17], xbs_fraction__54[18], xbs_fraction__54[19], xbs_fraction__54[20], xbs_fraction__54[21], xbs_fraction__54[22], xbs_fraction__54[23], xbs_fraction__54[24], xbs_fraction__54[25], xbs_fraction__54[26], xbs_fraction__54[27]};
  assign one_hot_171021 = {reverse_171013[27:0] == 28'h000_0000, reverse_171013[27] && reverse_171013[26:0] == 27'h000_0000, reverse_171013[26] && reverse_171013[25:0] == 26'h000_0000, reverse_171013[25] && reverse_171013[24:0] == 25'h000_0000, reverse_171013[24] && reverse_171013[23:0] == 24'h00_0000, reverse_171013[23] && reverse_171013[22:0] == 23'h00_0000, reverse_171013[22] && reverse_171013[21:0] == 22'h00_0000, reverse_171013[21] && reverse_171013[20:0] == 21'h00_0000, reverse_171013[20] && reverse_171013[19:0] == 20'h0_0000, reverse_171013[19] && reverse_171013[18:0] == 19'h0_0000, reverse_171013[18] && reverse_171013[17:0] == 18'h0_0000, reverse_171013[17] && reverse_171013[16:0] == 17'h0_0000, reverse_171013[16] && reverse_171013[15:0] == 16'h0000, reverse_171013[15] && reverse_171013[14:0] == 15'h0000, reverse_171013[14] && reverse_171013[13:0] == 14'h0000, reverse_171013[13] && reverse_171013[12:0] == 13'h0000, reverse_171013[12] && reverse_171013[11:0] == 12'h000, reverse_171013[11] && reverse_171013[10:0] == 11'h000, reverse_171013[10] && reverse_171013[9:0] == 10'h000, reverse_171013[9] && reverse_171013[8:0] == 9'h000, reverse_171013[8] && reverse_171013[7:0] == 8'h00, reverse_171013[7] && reverse_171013[6:0] == 7'h00, reverse_171013[6] && reverse_171013[5:0] == 6'h00, reverse_171013[5] && reverse_171013[4:0] == 5'h00, reverse_171013[4] && reverse_171013[3:0] == 4'h0, reverse_171013[3] && reverse_171013[2:0] == 3'h0, reverse_171013[2] && reverse_171013[1:0] == 2'h0, reverse_171013[1] && !reverse_171013[0], reverse_171013[0]};
  assign reverse_171022 = {xbs_fraction__72[0], xbs_fraction__72[1], xbs_fraction__72[2], xbs_fraction__72[3], xbs_fraction__72[4], xbs_fraction__72[5], xbs_fraction__72[6], xbs_fraction__72[7], xbs_fraction__72[8], xbs_fraction__72[9], xbs_fraction__72[10], xbs_fraction__72[11], xbs_fraction__72[12], xbs_fraction__72[13], xbs_fraction__72[14], xbs_fraction__72[15], xbs_fraction__72[16], xbs_fraction__72[17], xbs_fraction__72[18], xbs_fraction__72[19], xbs_fraction__72[20], xbs_fraction__72[21], xbs_fraction__72[22], xbs_fraction__72[23], xbs_fraction__72[24], xbs_fraction__72[25], xbs_fraction__72[26], xbs_fraction__72[27]};
  assign one_hot_171023 = {reverse_171015[27:0] == 28'h000_0000, reverse_171015[27] && reverse_171015[26:0] == 27'h000_0000, reverse_171015[26] && reverse_171015[25:0] == 26'h000_0000, reverse_171015[25] && reverse_171015[24:0] == 25'h000_0000, reverse_171015[24] && reverse_171015[23:0] == 24'h00_0000, reverse_171015[23] && reverse_171015[22:0] == 23'h00_0000, reverse_171015[22] && reverse_171015[21:0] == 22'h00_0000, reverse_171015[21] && reverse_171015[20:0] == 21'h00_0000, reverse_171015[20] && reverse_171015[19:0] == 20'h0_0000, reverse_171015[19] && reverse_171015[18:0] == 19'h0_0000, reverse_171015[18] && reverse_171015[17:0] == 18'h0_0000, reverse_171015[17] && reverse_171015[16:0] == 17'h0_0000, reverse_171015[16] && reverse_171015[15:0] == 16'h0000, reverse_171015[15] && reverse_171015[14:0] == 15'h0000, reverse_171015[14] && reverse_171015[13:0] == 14'h0000, reverse_171015[13] && reverse_171015[12:0] == 13'h0000, reverse_171015[12] && reverse_171015[11:0] == 12'h000, reverse_171015[11] && reverse_171015[10:0] == 11'h000, reverse_171015[10] && reverse_171015[9:0] == 10'h000, reverse_171015[9] && reverse_171015[8:0] == 9'h000, reverse_171015[8] && reverse_171015[7:0] == 8'h00, reverse_171015[7] && reverse_171015[6:0] == 7'h00, reverse_171015[6] && reverse_171015[5:0] == 6'h00, reverse_171015[5] && reverse_171015[4:0] == 5'h00, reverse_171015[4] && reverse_171015[3:0] == 4'h0, reverse_171015[3] && reverse_171015[2:0] == 3'h0, reverse_171015[2] && reverse_171015[1:0] == 2'h0, reverse_171015[1] && !reverse_171015[0], reverse_171015[0]};
  assign one_hot_171024 = {reverse_171016[27:0] == 28'h000_0000, reverse_171016[27] && reverse_171016[26:0] == 27'h000_0000, reverse_171016[26] && reverse_171016[25:0] == 26'h000_0000, reverse_171016[25] && reverse_171016[24:0] == 25'h000_0000, reverse_171016[24] && reverse_171016[23:0] == 24'h00_0000, reverse_171016[23] && reverse_171016[22:0] == 23'h00_0000, reverse_171016[22] && reverse_171016[21:0] == 22'h00_0000, reverse_171016[21] && reverse_171016[20:0] == 21'h00_0000, reverse_171016[20] && reverse_171016[19:0] == 20'h0_0000, reverse_171016[19] && reverse_171016[18:0] == 19'h0_0000, reverse_171016[18] && reverse_171016[17:0] == 18'h0_0000, reverse_171016[17] && reverse_171016[16:0] == 17'h0_0000, reverse_171016[16] && reverse_171016[15:0] == 16'h0000, reverse_171016[15] && reverse_171016[14:0] == 15'h0000, reverse_171016[14] && reverse_171016[13:0] == 14'h0000, reverse_171016[13] && reverse_171016[12:0] == 13'h0000, reverse_171016[12] && reverse_171016[11:0] == 12'h000, reverse_171016[11] && reverse_171016[10:0] == 11'h000, reverse_171016[10] && reverse_171016[9:0] == 10'h000, reverse_171016[9] && reverse_171016[8:0] == 9'h000, reverse_171016[8] && reverse_171016[7:0] == 8'h00, reverse_171016[7] && reverse_171016[6:0] == 7'h00, reverse_171016[6] && reverse_171016[5:0] == 6'h00, reverse_171016[5] && reverse_171016[4:0] == 5'h00, reverse_171016[4] && reverse_171016[3:0] == 4'h0, reverse_171016[3] && reverse_171016[2:0] == 3'h0, reverse_171016[2] && reverse_171016[1:0] == 2'h0, reverse_171016[1] && !reverse_171016[0], reverse_171016[0]};
  assign encode_171025 = {one_hot_171017[16] | one_hot_171017[17] | one_hot_171017[18] | one_hot_171017[19] | one_hot_171017[20] | one_hot_171017[21] | one_hot_171017[22] | one_hot_171017[23] | one_hot_171017[24] | one_hot_171017[25] | one_hot_171017[26] | one_hot_171017[27] | one_hot_171017[28], one_hot_171017[8] | one_hot_171017[9] | one_hot_171017[10] | one_hot_171017[11] | one_hot_171017[12] | one_hot_171017[13] | one_hot_171017[14] | one_hot_171017[15] | one_hot_171017[24] | one_hot_171017[25] | one_hot_171017[26] | one_hot_171017[27] | one_hot_171017[28], one_hot_171017[4] | one_hot_171017[5] | one_hot_171017[6] | one_hot_171017[7] | one_hot_171017[12] | one_hot_171017[13] | one_hot_171017[14] | one_hot_171017[15] | one_hot_171017[20] | one_hot_171017[21] | one_hot_171017[22] | one_hot_171017[23] | one_hot_171017[28], one_hot_171017[2] | one_hot_171017[3] | one_hot_171017[6] | one_hot_171017[7] | one_hot_171017[10] | one_hot_171017[11] | one_hot_171017[14] | one_hot_171017[15] | one_hot_171017[18] | one_hot_171017[19] | one_hot_171017[22] | one_hot_171017[23] | one_hot_171017[26] | one_hot_171017[27], one_hot_171017[1] | one_hot_171017[3] | one_hot_171017[5] | one_hot_171017[7] | one_hot_171017[9] | one_hot_171017[11] | one_hot_171017[13] | one_hot_171017[15] | one_hot_171017[17] | one_hot_171017[19] | one_hot_171017[21] | one_hot_171017[23] | one_hot_171017[25] | one_hot_171017[27]};
  assign one_hot_171026 = {reverse_171018[27:0] == 28'h000_0000, reverse_171018[27] && reverse_171018[26:0] == 27'h000_0000, reverse_171018[26] && reverse_171018[25:0] == 26'h000_0000, reverse_171018[25] && reverse_171018[24:0] == 25'h000_0000, reverse_171018[24] && reverse_171018[23:0] == 24'h00_0000, reverse_171018[23] && reverse_171018[22:0] == 23'h00_0000, reverse_171018[22] && reverse_171018[21:0] == 22'h00_0000, reverse_171018[21] && reverse_171018[20:0] == 21'h00_0000, reverse_171018[20] && reverse_171018[19:0] == 20'h0_0000, reverse_171018[19] && reverse_171018[18:0] == 19'h0_0000, reverse_171018[18] && reverse_171018[17:0] == 18'h0_0000, reverse_171018[17] && reverse_171018[16:0] == 17'h0_0000, reverse_171018[16] && reverse_171018[15:0] == 16'h0000, reverse_171018[15] && reverse_171018[14:0] == 15'h0000, reverse_171018[14] && reverse_171018[13:0] == 14'h0000, reverse_171018[13] && reverse_171018[12:0] == 13'h0000, reverse_171018[12] && reverse_171018[11:0] == 12'h000, reverse_171018[11] && reverse_171018[10:0] == 11'h000, reverse_171018[10] && reverse_171018[9:0] == 10'h000, reverse_171018[9] && reverse_171018[8:0] == 9'h000, reverse_171018[8] && reverse_171018[7:0] == 8'h00, reverse_171018[7] && reverse_171018[6:0] == 7'h00, reverse_171018[6] && reverse_171018[5:0] == 6'h00, reverse_171018[5] && reverse_171018[4:0] == 5'h00, reverse_171018[4] && reverse_171018[3:0] == 4'h0, reverse_171018[3] && reverse_171018[2:0] == 3'h0, reverse_171018[2] && reverse_171018[1:0] == 2'h0, reverse_171018[1] && !reverse_171018[0], reverse_171018[0]};
  assign encode_171027 = {one_hot_171019[16] | one_hot_171019[17] | one_hot_171019[18] | one_hot_171019[19] | one_hot_171019[20] | one_hot_171019[21] | one_hot_171019[22] | one_hot_171019[23] | one_hot_171019[24] | one_hot_171019[25] | one_hot_171019[26] | one_hot_171019[27] | one_hot_171019[28], one_hot_171019[8] | one_hot_171019[9] | one_hot_171019[10] | one_hot_171019[11] | one_hot_171019[12] | one_hot_171019[13] | one_hot_171019[14] | one_hot_171019[15] | one_hot_171019[24] | one_hot_171019[25] | one_hot_171019[26] | one_hot_171019[27] | one_hot_171019[28], one_hot_171019[4] | one_hot_171019[5] | one_hot_171019[6] | one_hot_171019[7] | one_hot_171019[12] | one_hot_171019[13] | one_hot_171019[14] | one_hot_171019[15] | one_hot_171019[20] | one_hot_171019[21] | one_hot_171019[22] | one_hot_171019[23] | one_hot_171019[28], one_hot_171019[2] | one_hot_171019[3] | one_hot_171019[6] | one_hot_171019[7] | one_hot_171019[10] | one_hot_171019[11] | one_hot_171019[14] | one_hot_171019[15] | one_hot_171019[18] | one_hot_171019[19] | one_hot_171019[22] | one_hot_171019[23] | one_hot_171019[26] | one_hot_171019[27], one_hot_171019[1] | one_hot_171019[3] | one_hot_171019[5] | one_hot_171019[7] | one_hot_171019[9] | one_hot_171019[11] | one_hot_171019[13] | one_hot_171019[15] | one_hot_171019[17] | one_hot_171019[19] | one_hot_171019[21] | one_hot_171019[23] | one_hot_171019[25] | one_hot_171019[27]};
  assign one_hot_171028 = {reverse_171020[27:0] == 28'h000_0000, reverse_171020[27] && reverse_171020[26:0] == 27'h000_0000, reverse_171020[26] && reverse_171020[25:0] == 26'h000_0000, reverse_171020[25] && reverse_171020[24:0] == 25'h000_0000, reverse_171020[24] && reverse_171020[23:0] == 24'h00_0000, reverse_171020[23] && reverse_171020[22:0] == 23'h00_0000, reverse_171020[22] && reverse_171020[21:0] == 22'h00_0000, reverse_171020[21] && reverse_171020[20:0] == 21'h00_0000, reverse_171020[20] && reverse_171020[19:0] == 20'h0_0000, reverse_171020[19] && reverse_171020[18:0] == 19'h0_0000, reverse_171020[18] && reverse_171020[17:0] == 18'h0_0000, reverse_171020[17] && reverse_171020[16:0] == 17'h0_0000, reverse_171020[16] && reverse_171020[15:0] == 16'h0000, reverse_171020[15] && reverse_171020[14:0] == 15'h0000, reverse_171020[14] && reverse_171020[13:0] == 14'h0000, reverse_171020[13] && reverse_171020[12:0] == 13'h0000, reverse_171020[12] && reverse_171020[11:0] == 12'h000, reverse_171020[11] && reverse_171020[10:0] == 11'h000, reverse_171020[10] && reverse_171020[9:0] == 10'h000, reverse_171020[9] && reverse_171020[8:0] == 9'h000, reverse_171020[8] && reverse_171020[7:0] == 8'h00, reverse_171020[7] && reverse_171020[6:0] == 7'h00, reverse_171020[6] && reverse_171020[5:0] == 6'h00, reverse_171020[5] && reverse_171020[4:0] == 5'h00, reverse_171020[4] && reverse_171020[3:0] == 4'h0, reverse_171020[3] && reverse_171020[2:0] == 3'h0, reverse_171020[2] && reverse_171020[1:0] == 2'h0, reverse_171020[1] && !reverse_171020[0], reverse_171020[0]};
  assign encode_171029 = {one_hot_171021[16] | one_hot_171021[17] | one_hot_171021[18] | one_hot_171021[19] | one_hot_171021[20] | one_hot_171021[21] | one_hot_171021[22] | one_hot_171021[23] | one_hot_171021[24] | one_hot_171021[25] | one_hot_171021[26] | one_hot_171021[27] | one_hot_171021[28], one_hot_171021[8] | one_hot_171021[9] | one_hot_171021[10] | one_hot_171021[11] | one_hot_171021[12] | one_hot_171021[13] | one_hot_171021[14] | one_hot_171021[15] | one_hot_171021[24] | one_hot_171021[25] | one_hot_171021[26] | one_hot_171021[27] | one_hot_171021[28], one_hot_171021[4] | one_hot_171021[5] | one_hot_171021[6] | one_hot_171021[7] | one_hot_171021[12] | one_hot_171021[13] | one_hot_171021[14] | one_hot_171021[15] | one_hot_171021[20] | one_hot_171021[21] | one_hot_171021[22] | one_hot_171021[23] | one_hot_171021[28], one_hot_171021[2] | one_hot_171021[3] | one_hot_171021[6] | one_hot_171021[7] | one_hot_171021[10] | one_hot_171021[11] | one_hot_171021[14] | one_hot_171021[15] | one_hot_171021[18] | one_hot_171021[19] | one_hot_171021[22] | one_hot_171021[23] | one_hot_171021[26] | one_hot_171021[27], one_hot_171021[1] | one_hot_171021[3] | one_hot_171021[5] | one_hot_171021[7] | one_hot_171021[9] | one_hot_171021[11] | one_hot_171021[13] | one_hot_171021[15] | one_hot_171021[17] | one_hot_171021[19] | one_hot_171021[21] | one_hot_171021[23] | one_hot_171021[25] | one_hot_171021[27]};
  assign one_hot_171030 = {reverse_171022[27:0] == 28'h000_0000, reverse_171022[27] && reverse_171022[26:0] == 27'h000_0000, reverse_171022[26] && reverse_171022[25:0] == 26'h000_0000, reverse_171022[25] && reverse_171022[24:0] == 25'h000_0000, reverse_171022[24] && reverse_171022[23:0] == 24'h00_0000, reverse_171022[23] && reverse_171022[22:0] == 23'h00_0000, reverse_171022[22] && reverse_171022[21:0] == 22'h00_0000, reverse_171022[21] && reverse_171022[20:0] == 21'h00_0000, reverse_171022[20] && reverse_171022[19:0] == 20'h0_0000, reverse_171022[19] && reverse_171022[18:0] == 19'h0_0000, reverse_171022[18] && reverse_171022[17:0] == 18'h0_0000, reverse_171022[17] && reverse_171022[16:0] == 17'h0_0000, reverse_171022[16] && reverse_171022[15:0] == 16'h0000, reverse_171022[15] && reverse_171022[14:0] == 15'h0000, reverse_171022[14] && reverse_171022[13:0] == 14'h0000, reverse_171022[13] && reverse_171022[12:0] == 13'h0000, reverse_171022[12] && reverse_171022[11:0] == 12'h000, reverse_171022[11] && reverse_171022[10:0] == 11'h000, reverse_171022[10] && reverse_171022[9:0] == 10'h000, reverse_171022[9] && reverse_171022[8:0] == 9'h000, reverse_171022[8] && reverse_171022[7:0] == 8'h00, reverse_171022[7] && reverse_171022[6:0] == 7'h00, reverse_171022[6] && reverse_171022[5:0] == 6'h00, reverse_171022[5] && reverse_171022[4:0] == 5'h00, reverse_171022[4] && reverse_171022[3:0] == 4'h0, reverse_171022[3] && reverse_171022[2:0] == 3'h0, reverse_171022[2] && reverse_171022[1:0] == 2'h0, reverse_171022[1] && !reverse_171022[0], reverse_171022[0]};
  assign encode_171031 = {one_hot_171023[16] | one_hot_171023[17] | one_hot_171023[18] | one_hot_171023[19] | one_hot_171023[20] | one_hot_171023[21] | one_hot_171023[22] | one_hot_171023[23] | one_hot_171023[24] | one_hot_171023[25] | one_hot_171023[26] | one_hot_171023[27] | one_hot_171023[28], one_hot_171023[8] | one_hot_171023[9] | one_hot_171023[10] | one_hot_171023[11] | one_hot_171023[12] | one_hot_171023[13] | one_hot_171023[14] | one_hot_171023[15] | one_hot_171023[24] | one_hot_171023[25] | one_hot_171023[26] | one_hot_171023[27] | one_hot_171023[28], one_hot_171023[4] | one_hot_171023[5] | one_hot_171023[6] | one_hot_171023[7] | one_hot_171023[12] | one_hot_171023[13] | one_hot_171023[14] | one_hot_171023[15] | one_hot_171023[20] | one_hot_171023[21] | one_hot_171023[22] | one_hot_171023[23] | one_hot_171023[28], one_hot_171023[2] | one_hot_171023[3] | one_hot_171023[6] | one_hot_171023[7] | one_hot_171023[10] | one_hot_171023[11] | one_hot_171023[14] | one_hot_171023[15] | one_hot_171023[18] | one_hot_171023[19] | one_hot_171023[22] | one_hot_171023[23] | one_hot_171023[26] | one_hot_171023[27], one_hot_171023[1] | one_hot_171023[3] | one_hot_171023[5] | one_hot_171023[7] | one_hot_171023[9] | one_hot_171023[11] | one_hot_171023[13] | one_hot_171023[15] | one_hot_171023[17] | one_hot_171023[19] | one_hot_171023[21] | one_hot_171023[23] | one_hot_171023[25] | one_hot_171023[27]};
  assign encode_171032 = {one_hot_171024[16] | one_hot_171024[17] | one_hot_171024[18] | one_hot_171024[19] | one_hot_171024[20] | one_hot_171024[21] | one_hot_171024[22] | one_hot_171024[23] | one_hot_171024[24] | one_hot_171024[25] | one_hot_171024[26] | one_hot_171024[27] | one_hot_171024[28], one_hot_171024[8] | one_hot_171024[9] | one_hot_171024[10] | one_hot_171024[11] | one_hot_171024[12] | one_hot_171024[13] | one_hot_171024[14] | one_hot_171024[15] | one_hot_171024[24] | one_hot_171024[25] | one_hot_171024[26] | one_hot_171024[27] | one_hot_171024[28], one_hot_171024[4] | one_hot_171024[5] | one_hot_171024[6] | one_hot_171024[7] | one_hot_171024[12] | one_hot_171024[13] | one_hot_171024[14] | one_hot_171024[15] | one_hot_171024[20] | one_hot_171024[21] | one_hot_171024[22] | one_hot_171024[23] | one_hot_171024[28], one_hot_171024[2] | one_hot_171024[3] | one_hot_171024[6] | one_hot_171024[7] | one_hot_171024[10] | one_hot_171024[11] | one_hot_171024[14] | one_hot_171024[15] | one_hot_171024[18] | one_hot_171024[19] | one_hot_171024[22] | one_hot_171024[23] | one_hot_171024[26] | one_hot_171024[27], one_hot_171024[1] | one_hot_171024[3] | one_hot_171024[5] | one_hot_171024[7] | one_hot_171024[9] | one_hot_171024[11] | one_hot_171024[13] | one_hot_171024[15] | one_hot_171024[17] | one_hot_171024[19] | one_hot_171024[21] | one_hot_171024[23] | one_hot_171024[25] | one_hot_171024[27]};
  assign encode_171034 = {one_hot_171026[16] | one_hot_171026[17] | one_hot_171026[18] | one_hot_171026[19] | one_hot_171026[20] | one_hot_171026[21] | one_hot_171026[22] | one_hot_171026[23] | one_hot_171026[24] | one_hot_171026[25] | one_hot_171026[26] | one_hot_171026[27] | one_hot_171026[28], one_hot_171026[8] | one_hot_171026[9] | one_hot_171026[10] | one_hot_171026[11] | one_hot_171026[12] | one_hot_171026[13] | one_hot_171026[14] | one_hot_171026[15] | one_hot_171026[24] | one_hot_171026[25] | one_hot_171026[26] | one_hot_171026[27] | one_hot_171026[28], one_hot_171026[4] | one_hot_171026[5] | one_hot_171026[6] | one_hot_171026[7] | one_hot_171026[12] | one_hot_171026[13] | one_hot_171026[14] | one_hot_171026[15] | one_hot_171026[20] | one_hot_171026[21] | one_hot_171026[22] | one_hot_171026[23] | one_hot_171026[28], one_hot_171026[2] | one_hot_171026[3] | one_hot_171026[6] | one_hot_171026[7] | one_hot_171026[10] | one_hot_171026[11] | one_hot_171026[14] | one_hot_171026[15] | one_hot_171026[18] | one_hot_171026[19] | one_hot_171026[22] | one_hot_171026[23] | one_hot_171026[26] | one_hot_171026[27], one_hot_171026[1] | one_hot_171026[3] | one_hot_171026[5] | one_hot_171026[7] | one_hot_171026[9] | one_hot_171026[11] | one_hot_171026[13] | one_hot_171026[15] | one_hot_171026[17] | one_hot_171026[19] | one_hot_171026[21] | one_hot_171026[23] | one_hot_171026[25] | one_hot_171026[27]};
  assign encode_171036 = {one_hot_171028[16] | one_hot_171028[17] | one_hot_171028[18] | one_hot_171028[19] | one_hot_171028[20] | one_hot_171028[21] | one_hot_171028[22] | one_hot_171028[23] | one_hot_171028[24] | one_hot_171028[25] | one_hot_171028[26] | one_hot_171028[27] | one_hot_171028[28], one_hot_171028[8] | one_hot_171028[9] | one_hot_171028[10] | one_hot_171028[11] | one_hot_171028[12] | one_hot_171028[13] | one_hot_171028[14] | one_hot_171028[15] | one_hot_171028[24] | one_hot_171028[25] | one_hot_171028[26] | one_hot_171028[27] | one_hot_171028[28], one_hot_171028[4] | one_hot_171028[5] | one_hot_171028[6] | one_hot_171028[7] | one_hot_171028[12] | one_hot_171028[13] | one_hot_171028[14] | one_hot_171028[15] | one_hot_171028[20] | one_hot_171028[21] | one_hot_171028[22] | one_hot_171028[23] | one_hot_171028[28], one_hot_171028[2] | one_hot_171028[3] | one_hot_171028[6] | one_hot_171028[7] | one_hot_171028[10] | one_hot_171028[11] | one_hot_171028[14] | one_hot_171028[15] | one_hot_171028[18] | one_hot_171028[19] | one_hot_171028[22] | one_hot_171028[23] | one_hot_171028[26] | one_hot_171028[27], one_hot_171028[1] | one_hot_171028[3] | one_hot_171028[5] | one_hot_171028[7] | one_hot_171028[9] | one_hot_171028[11] | one_hot_171028[13] | one_hot_171028[15] | one_hot_171028[17] | one_hot_171028[19] | one_hot_171028[21] | one_hot_171028[23] | one_hot_171028[25] | one_hot_171028[27]};
  assign encode_171038 = {one_hot_171030[16] | one_hot_171030[17] | one_hot_171030[18] | one_hot_171030[19] | one_hot_171030[20] | one_hot_171030[21] | one_hot_171030[22] | one_hot_171030[23] | one_hot_171030[24] | one_hot_171030[25] | one_hot_171030[26] | one_hot_171030[27] | one_hot_171030[28], one_hot_171030[8] | one_hot_171030[9] | one_hot_171030[10] | one_hot_171030[11] | one_hot_171030[12] | one_hot_171030[13] | one_hot_171030[14] | one_hot_171030[15] | one_hot_171030[24] | one_hot_171030[25] | one_hot_171030[26] | one_hot_171030[27] | one_hot_171030[28], one_hot_171030[4] | one_hot_171030[5] | one_hot_171030[6] | one_hot_171030[7] | one_hot_171030[12] | one_hot_171030[13] | one_hot_171030[14] | one_hot_171030[15] | one_hot_171030[20] | one_hot_171030[21] | one_hot_171030[22] | one_hot_171030[23] | one_hot_171030[28], one_hot_171030[2] | one_hot_171030[3] | one_hot_171030[6] | one_hot_171030[7] | one_hot_171030[10] | one_hot_171030[11] | one_hot_171030[14] | one_hot_171030[15] | one_hot_171030[18] | one_hot_171030[19] | one_hot_171030[22] | one_hot_171030[23] | one_hot_171030[26] | one_hot_171030[27], one_hot_171030[1] | one_hot_171030[3] | one_hot_171030[5] | one_hot_171030[7] | one_hot_171030[9] | one_hot_171030[11] | one_hot_171030[13] | one_hot_171030[15] | one_hot_171030[17] | one_hot_171030[19] | one_hot_171030[21] | one_hot_171030[23] | one_hot_171030[25] | one_hot_171030[27]};
  assign cancel__18 = |encode_171025[4:1];
  assign carry_bit__17 = xbs_fraction__17[27];
  assign result_fraction__526 = 23'h00_0000;
  assign cancel__36 = |encode_171027[4:1];
  assign carry_bit__36 = xbs_fraction__35[27];
  assign result_fraction__593 = 23'h00_0000;
  assign cancel__55 = |encode_171029[4:1];
  assign carry_bit__55 = xbs_fraction__53[27];
  assign result_fraction__660 = 23'h00_0000;
  assign cancel__74 = |encode_171031[4:1];
  assign carry_bit__74 = xbs_fraction__71[27];
  assign result_fraction__739 = 23'h00_0000;
  assign cancel__9 = |encode_171032[4:1];
  assign carry_bit__18 = xbs_fraction__18[27];
  assign result_fraction__527 = 23'h00_0000;
  assign leading_zeroes__17 = {result_fraction__526, encode_171025};
  assign cancel__37 = |encode_171034[4:1];
  assign carry_bit__37 = xbs_fraction__36[27];
  assign result_fraction__594 = 23'h00_0000;
  assign leading_zeroes__36 = {result_fraction__593, encode_171027};
  assign cancel__56 = |encode_171036[4:1];
  assign carry_bit__56 = xbs_fraction__54[27];
  assign result_fraction__661 = 23'h00_0000;
  assign leading_zeroes__55 = {result_fraction__660, encode_171029};
  assign cancel__75 = |encode_171038[4:1];
  assign carry_bit__75 = xbs_fraction__72[27];
  assign result_fraction__740 = 23'h00_0000;
  assign leading_zeroes__74 = {result_fraction__739, encode_171031};
  assign leading_zeroes__18 = {result_fraction__527, encode_171032};
  assign carry_fraction__34 = xbs_fraction__17[27:1];
  assign add_171104 = leading_zeroes__17 + 28'hfff_ffff;
  assign leading_zeroes__37 = {result_fraction__594, encode_171034};
  assign carry_fraction__71 = xbs_fraction__35[27:1];
  assign add_171117 = leading_zeroes__36 + 28'hfff_ffff;
  assign leading_zeroes__56 = {result_fraction__661, encode_171036};
  assign carry_fraction__109 = xbs_fraction__53[27:1];
  assign add_171130 = leading_zeroes__55 + 28'hfff_ffff;
  assign leading_zeroes__75 = {result_fraction__740, encode_171038};
  assign carry_fraction__147 = xbs_fraction__71[27:1];
  assign add_171143 = leading_zeroes__74 + 28'hfff_ffff;
  assign carry_fraction__17 = xbs_fraction__18[27:1];
  assign add_171150 = leading_zeroes__18 + 28'hfff_ffff;
  assign concat_171151 = {~(carry_bit__17 | cancel__18), ~(carry_bit__17 | ~cancel__18), ~(~carry_bit__17 | cancel__18)};
  assign carry_fraction__35 = carry_fraction__34 | {26'h000_0000, xbs_fraction__17[0]};
  assign cancel_fraction__17 = add_171104 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__17[26:0] << add_171104;
  assign carry_fraction__72 = xbs_fraction__36[27:1];
  assign add_171160 = leading_zeroes__37 + 28'hfff_ffff;
  assign concat_171161 = {~(carry_bit__36 | cancel__36), ~(carry_bit__36 | ~cancel__36), ~(~carry_bit__36 | cancel__36)};
  assign carry_fraction__73 = carry_fraction__71 | {26'h000_0000, xbs_fraction__35[0]};
  assign cancel_fraction__36 = add_171117 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__35[26:0] << add_171117;
  assign carry_fraction__110 = xbs_fraction__54[27:1];
  assign add_171170 = leading_zeroes__56 + 28'hfff_ffff;
  assign concat_171171 = {~(carry_bit__55 | cancel__55), ~(carry_bit__55 | ~cancel__55), ~(~carry_bit__55 | cancel__55)};
  assign carry_fraction__111 = carry_fraction__109 | {26'h000_0000, xbs_fraction__53[0]};
  assign cancel_fraction__55 = add_171130 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__53[26:0] << add_171130;
  assign carry_fraction__148 = xbs_fraction__72[27:1];
  assign add_171180 = leading_zeroes__75 + 28'hfff_ffff;
  assign concat_171181 = {~(carry_bit__74 | cancel__74), ~(carry_bit__74 | ~cancel__74), ~(~carry_bit__74 | cancel__74)};
  assign carry_fraction__149 = carry_fraction__147 | {26'h000_0000, xbs_fraction__71[0]};
  assign cancel_fraction__74 = add_171143 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__71[26:0] << add_171143;
  assign concat_171184 = {~(carry_bit__18 | cancel__9), ~(carry_bit__18 | ~cancel__9), ~(~carry_bit__18 | cancel__9)};
  assign carry_fraction__36 = carry_fraction__17 | {26'h000_0000, xbs_fraction__18[0]};
  assign cancel_fraction__18 = add_171150 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__18[26:0] << add_171150;
  assign shifted_fraction__17 = carry_fraction__35 & {27{concat_171151[0]}} | cancel_fraction__17 & {27{concat_171151[1]}} | xbs_fraction__17[26:0] & {27{concat_171151[2]}};
  assign concat_171188 = {~(carry_bit__37 | cancel__37), ~(carry_bit__37 | ~cancel__37), ~(~carry_bit__37 | cancel__37)};
  assign carry_fraction__74 = carry_fraction__72 | {26'h000_0000, xbs_fraction__36[0]};
  assign cancel_fraction__37 = add_171160 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__36[26:0] << add_171160;
  assign shifted_fraction__36 = carry_fraction__73 & {27{concat_171161[0]}} | cancel_fraction__36 & {27{concat_171161[1]}} | xbs_fraction__35[26:0] & {27{concat_171161[2]}};
  assign concat_171192 = {~(carry_bit__56 | cancel__56), ~(carry_bit__56 | ~cancel__56), ~(~carry_bit__56 | cancel__56)};
  assign carry_fraction__112 = carry_fraction__110 | {26'h000_0000, xbs_fraction__54[0]};
  assign cancel_fraction__56 = add_171170 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__54[26:0] << add_171170;
  assign shifted_fraction__55 = carry_fraction__111 & {27{concat_171171[0]}} | cancel_fraction__55 & {27{concat_171171[1]}} | xbs_fraction__53[26:0] & {27{concat_171171[2]}};
  assign concat_171196 = {~(carry_bit__75 | cancel__75), ~(carry_bit__75 | ~cancel__75), ~(~carry_bit__75 | cancel__75)};
  assign carry_fraction__150 = carry_fraction__148 | {26'h000_0000, xbs_fraction__72[0]};
  assign cancel_fraction__75 = add_171180 >= 28'h000_001b ? 27'h000_0000 : xbs_fraction__72[26:0] << add_171180;
  assign shifted_fraction__74 = carry_fraction__149 & {27{concat_171181[0]}} | cancel_fraction__74 & {27{concat_171181[1]}} | xbs_fraction__71[26:0] & {27{concat_171181[2]}};
  assign shifted_fraction__18 = carry_fraction__36 & {27{concat_171184[0]}} | cancel_fraction__18 & {27{concat_171184[1]}} | xbs_fraction__18[26:0] & {27{concat_171184[2]}};
  assign result_sign__1092 = 1'h0;
  assign shifted_fraction__37 = carry_fraction__74 & {27{concat_171188[0]}} | cancel_fraction__37 & {27{concat_171188[1]}} | xbs_fraction__36[26:0] & {27{concat_171188[2]}};
  assign result_sign__1093 = 1'h0;
  assign shifted_fraction__56 = carry_fraction__112 & {27{concat_171192[0]}} | cancel_fraction__56 & {27{concat_171192[1]}} | xbs_fraction__54[26:0] & {27{concat_171192[2]}};
  assign result_sign__1094 = 1'h0;
  assign shifted_fraction__75 = carry_fraction__150 & {27{concat_171196[0]}} | cancel_fraction__75 & {27{concat_171196[1]}} | xbs_fraction__72[26:0] & {27{concat_171196[2]}};
  assign result_sign__1095 = 1'h0;
  assign result_sign__1096 = 1'h0;
  assign normal_chunk__17 = shifted_fraction__17[2:0];
  assign fraction_shift__257 = 3'h4;
  assign half_way_chunk__17 = shifted_fraction__17[3:2];
  assign result_sign__1097 = 1'h0;
  assign normal_chunk__36 = shifted_fraction__36[2:0];
  assign fraction_shift__292 = 3'h4;
  assign half_way_chunk__36 = shifted_fraction__36[3:2];
  assign result_sign__1098 = 1'h0;
  assign normal_chunk__55 = shifted_fraction__55[2:0];
  assign fraction_shift__327 = 3'h4;
  assign half_way_chunk__55 = shifted_fraction__55[3:2];
  assign result_sign__1099 = 1'h0;
  assign normal_chunk__74 = shifted_fraction__74[2:0];
  assign fraction_shift__362 = 3'h4;
  assign half_way_chunk__74 = shifted_fraction__74[3:2];
  assign normal_chunk__18 = shifted_fraction__18[2:0];
  assign fraction_shift__258 = 3'h4;
  assign half_way_chunk__18 = shifted_fraction__18[3:2];
  assign result_sign__460 = 1'h0;
  assign add_171253 = {result_sign__1092, shifted_fraction__17[26:3]} + 25'h000_0001;
  assign normal_chunk__37 = shifted_fraction__37[2:0];
  assign fraction_shift__293 = 3'h4;
  assign half_way_chunk__37 = shifted_fraction__37[3:2];
  assign result_sign__557 = 1'h0;
  assign add_171263 = {result_sign__1093, shifted_fraction__36[26:3]} + 25'h000_0001;
  assign normal_chunk__56 = shifted_fraction__56[2:0];
  assign fraction_shift__328 = 3'h4;
  assign half_way_chunk__56 = shifted_fraction__56[3:2];
  assign result_sign__659 = 1'h0;
  assign add_171273 = {result_sign__1094, shifted_fraction__55[26:3]} + 25'h000_0001;
  assign normal_chunk__75 = shifted_fraction__75[2:0];
  assign fraction_shift__363 = 3'h4;
  assign half_way_chunk__75 = shifted_fraction__75[3:2];
  assign result_sign__771 = 1'h0;
  assign add_171283 = {result_sign__1095, shifted_fraction__74[26:3]} + 25'h000_0001;
  assign result_sign__461 = 1'h0;
  assign add_171287 = {result_sign__1096, shifted_fraction__18[26:3]} + 25'h000_0001;
  assign do_round_up__35 = normal_chunk__17 > fraction_shift__257 | half_way_chunk__17 == 2'h3;
  assign result_sign__558 = 1'h0;
  assign add_171294 = {result_sign__1097, shifted_fraction__37[26:3]} + 25'h000_0001;
  assign do_round_up__74 = normal_chunk__36 > fraction_shift__292 | half_way_chunk__36 == 2'h3;
  assign result_sign__660 = 1'h0;
  assign add_171301 = {result_sign__1098, shifted_fraction__56[26:3]} + 25'h000_0001;
  assign do_round_up__113 = normal_chunk__55 > fraction_shift__327 | half_way_chunk__55 == 2'h3;
  assign result_sign__772 = 1'h0;
  assign add_171308 = {result_sign__1099, shifted_fraction__75[26:3]} + 25'h000_0001;
  assign do_round_up__152 = normal_chunk__74 > fraction_shift__362 | half_way_chunk__74 == 2'h3;
  assign do_round_up__36 = normal_chunk__18 > fraction_shift__258 | half_way_chunk__18 == 2'h3;
  assign rounded_fraction__17 = do_round_up__35 ? {add_171253, normal_chunk__17} : {result_sign__460, shifted_fraction__17};
  assign do_round_up__75 = normal_chunk__37 > fraction_shift__293 | half_way_chunk__37 == 2'h3;
  assign rounded_fraction__36 = do_round_up__74 ? {add_171263, normal_chunk__36} : {result_sign__557, shifted_fraction__36};
  assign do_round_up__114 = normal_chunk__56 > fraction_shift__328 | half_way_chunk__56 == 2'h3;
  assign rounded_fraction__55 = do_round_up__113 ? {add_171273, normal_chunk__55} : {result_sign__659, shifted_fraction__55};
  assign do_round_up__153 = normal_chunk__75 > fraction_shift__363 | half_way_chunk__75 == 2'h3;
  assign rounded_fraction__74 = do_round_up__152 ? {add_171283, normal_chunk__74} : {result_sign__771, shifted_fraction__74};
  assign rounded_fraction__18 = do_round_up__36 ? {add_171287, normal_chunk__18} : {result_sign__461, shifted_fraction__18};
  assign result_sign__462 = 1'h0;
  assign x_bexp__590 = 8'h00;
  assign rounding_carry__17 = rounded_fraction__17[27];
  assign rounded_fraction__37 = do_round_up__75 ? {add_171294, normal_chunk__37} : {result_sign__558, shifted_fraction__37};
  assign result_sign__559 = 1'h0;
  assign x_bexp__608 = 8'h00;
  assign rounding_carry__36 = rounded_fraction__36[27];
  assign rounded_fraction__56 = do_round_up__114 ? {add_171301, normal_chunk__56} : {result_sign__660, shifted_fraction__56};
  assign result_sign__661 = 1'h0;
  assign x_bexp__626 = 8'h00;
  assign rounding_carry__55 = rounded_fraction__55[27];
  assign rounded_fraction__75 = do_round_up__153 ? {add_171308, normal_chunk__75} : {result_sign__772, shifted_fraction__75};
  assign result_sign__773 = 1'h0;
  assign x_bexp__644 = 8'h00;
  assign rounding_carry__74 = rounded_fraction__74[27];
  assign result_sign__463 = 1'h0;
  assign x_bexp__591 = 8'h00;
  assign rounding_carry__18 = rounded_fraction__18[27];
  assign result_sign__560 = 1'h0;
  assign x_bexp__609 = 8'h00;
  assign rounding_carry__37 = rounded_fraction__37[27];
  assign result_sign__662 = 1'h0;
  assign x_bexp__627 = 8'h00;
  assign rounding_carry__56 = rounded_fraction__56[27];
  assign result_sign__774 = 1'h0;
  assign x_bexp__645 = 8'h00;
  assign rounding_carry__75 = rounded_fraction__75[27];
  assign result_sign__464 = 1'h0;
  assign add_171367 = {result_sign__462, x_bexp__142} + {x_bexp__590, rounding_carry__17};
  assign result_sign__561 = 1'h0;
  assign add_171373 = {result_sign__559, x_bexp__283} + {x_bexp__608, rounding_carry__36};
  assign result_sign__663 = 1'h0;
  assign add_171379 = {result_sign__661, x_bexp__427} + {x_bexp__626, rounding_carry__55};
  assign result_sign__775 = 1'h0;
  assign add_171385 = {result_sign__773, x_bexp__571} + {x_bexp__644, rounding_carry__74};
  assign result_sign__465 = 1'h0;
  assign add_171389 = {result_sign__463, x_bexp__70} + {x_bexp__591, rounding_carry__18};
  assign result_sign__562 = 1'h0;
  assign add_171398 = {result_sign__560, x_bexp__284} + {x_bexp__609, rounding_carry__37};
  assign result_sign__664 = 1'h0;
  assign add_171407 = {result_sign__662, x_bexp__428} + {x_bexp__627, rounding_carry__56};
  assign result_sign__776 = 1'h0;
  assign add_171416 = {result_sign__774, x_bexp__572} + {x_bexp__645, rounding_carry__75};
  assign add_171429 = {result_sign__464, add_171367} + 10'h001;
  assign add_171437 = {result_sign__561, add_171373} + 10'h001;
  assign add_171445 = {result_sign__663, add_171379} + 10'h001;
  assign add_171453 = {result_sign__775, add_171385} + 10'h001;
  assign add_171456 = {result_sign__465, add_171389} + 10'h001;
  assign wide_exponent__51 = add_171429 - {5'h00, encode_171025};
  assign add_171461 = {result_sign__562, add_171398} + 10'h001;
  assign wide_exponent__106 = add_171437 - {5'h00, encode_171027};
  assign add_171466 = {result_sign__664, add_171407} + 10'h001;
  assign wide_exponent__163 = add_171445 - {5'h00, encode_171029};
  assign add_171471 = {result_sign__776, add_171416} + 10'h001;
  assign wide_exponent__220 = add_171453 - {5'h00, encode_171031};
  assign wide_exponent__25 = add_171456 - {5'h00, encode_171032};
  assign wide_exponent__52 = wide_exponent__51 & {10{add_170950 != 26'h000_0000 | xddend_y__17[2:0] != 3'h0}};
  assign wide_exponent__107 = add_171461 - {5'h00, encode_171034};
  assign wide_exponent__108 = wide_exponent__106 & {10{add_170953 != 26'h000_0000 | xddend_y__35[2:0] != 3'h0}};
  assign wide_exponent__164 = add_171466 - {5'h00, encode_171036};
  assign wide_exponent__165 = wide_exponent__163 & {10{add_170956 != 26'h000_0000 | xddend_y__53[2:0] != 3'h0}};
  assign wide_exponent__221 = add_171471 - {5'h00, encode_171038};
  assign wide_exponent__222 = wide_exponent__220 & {10{add_170959 != 26'h000_0000 | xddend_y__71[2:0] != 3'h0}};
  assign wide_exponent__26 = wide_exponent__25 & {10{add_170960 != 26'h000_0000 | xddend_y__18[2:0] != 3'h0}};
  assign wide_exponent__109 = wide_exponent__107 & {10{add_170963 != 26'h000_0000 | xddend_y__36[2:0] != 3'h0}};
  assign wide_exponent__166 = wide_exponent__164 & {10{add_170966 != 26'h000_0000 | xddend_y__54[2:0] != 3'h0}};
  assign wide_exponent__223 = wide_exponent__221 & {10{add_170969 != 26'h000_0000 | xddend_y__72[2:0] != 3'h0}};
  assign high_exp__130 = 8'hff;
  assign result_fraction__528 = 23'h00_0000;
  assign high_exp__131 = 8'hff;
  assign result_fraction__529 = 23'h00_0000;
  assign wide_exponent__53 = wide_exponent__52[8:0] & {9{~wide_exponent__52[9]}};
  assign high_exp__195 = 8'hff;
  assign result_fraction__595 = 23'h00_0000;
  assign high_exp__196 = 8'hff;
  assign result_fraction__596 = 23'h00_0000;
  assign wide_exponent__110 = wide_exponent__108[8:0] & {9{~wide_exponent__108[9]}};
  assign high_exp__263 = 8'hff;
  assign result_fraction__662 = 23'h00_0000;
  assign high_exp__264 = 8'hff;
  assign result_fraction__663 = 23'h00_0000;
  assign wide_exponent__167 = wide_exponent__165[8:0] & {9{~wide_exponent__165[9]}};
  assign high_exp__337 = 8'hff;
  assign result_fraction__741 = 23'h00_0000;
  assign high_exp__338 = 8'hff;
  assign result_fraction__742 = 23'h00_0000;
  assign wide_exponent__224 = wide_exponent__222[8:0] & {9{~wide_exponent__222[9]}};
  assign high_exp__132 = 8'hff;
  assign result_fraction__530 = 23'h00_0000;
  assign high_exp__133 = 8'hff;
  assign result_fraction__531 = 23'h00_0000;
  assign wide_exponent__54 = wide_exponent__26[8:0] & {9{~wide_exponent__26[9]}};
  assign eq_171549 = x_bexp__142 == high_exp__130;
  assign eq_171550 = x_fraction__142 == result_fraction__528;
  assign eq_171551 = prod_bexp__70 == high_exp__131;
  assign eq_171552 = prod_fraction__51 == result_fraction__529;
  assign high_exp__381 = 8'hff;
  assign result_fraction__787 = 23'h00_0000;
  assign high_exp__382 = 8'hff;
  assign result_fraction__788 = 23'h00_0000;
  assign high_exp__197 = 8'hff;
  assign result_fraction__597 = 23'h00_0000;
  assign high_exp__198 = 8'hff;
  assign result_fraction__598 = 23'h00_0000;
  assign wide_exponent__111 = wide_exponent__109[8:0] & {9{~wide_exponent__109[9]}};
  assign eq_171563 = x_bexp__283 == high_exp__195;
  assign eq_171564 = x_fraction__283 == result_fraction__595;
  assign eq_171565 = prod_bexp__139 == high_exp__196;
  assign eq_171566 = prod_fraction__103 == result_fraction__596;
  assign high_exp__413 = 8'hff;
  assign result_fraction__820 = 23'h00_0000;
  assign high_exp__414 = 8'hff;
  assign result_fraction__821 = 23'h00_0000;
  assign high_exp__265 = 8'hff;
  assign result_fraction__664 = 23'h00_0000;
  assign high_exp__266 = 8'hff;
  assign result_fraction__665 = 23'h00_0000;
  assign wide_exponent__168 = wide_exponent__166[8:0] & {9{~wide_exponent__166[9]}};
  assign eq_171577 = x_bexp__427 == high_exp__263;
  assign eq_171578 = x_fraction__427 == result_fraction__662;
  assign eq_171579 = prod_bexp__211 == high_exp__264;
  assign eq_171580 = prod_fraction__157 == result_fraction__663;
  assign high_exp__445 = 8'hff;
  assign result_fraction__853 = 23'h00_0000;
  assign high_exp__446 = 8'hff;
  assign result_fraction__854 = 23'h00_0000;
  assign high_exp__339 = 8'hff;
  assign result_fraction__743 = 23'h00_0000;
  assign high_exp__340 = 8'hff;
  assign result_fraction__744 = 23'h00_0000;
  assign wide_exponent__225 = wide_exponent__223[8:0] & {9{~wide_exponent__223[9]}};
  assign eq_171591 = x_bexp__571 == high_exp__337;
  assign eq_171592 = x_fraction__571 == result_fraction__741;
  assign eq_171593 = prod_bexp__283 == high_exp__338;
  assign eq_171594 = prod_fraction__211 == result_fraction__742;
  assign high_exp__477 = 8'hff;
  assign result_fraction__886 = 23'h00_0000;
  assign high_exp__478 = 8'hff;
  assign result_fraction__887 = 23'h00_0000;
  assign eq_171600 = x_bexp__70 == high_exp__132;
  assign eq_171601 = x_fraction__70 == result_fraction__530;
  assign eq_171602 = prod_bexp__34 == high_exp__133;
  assign eq_171603 = prod_fraction__25 == result_fraction__531;
  assign high_exp__379 = 8'hff;
  assign result_fraction__785 = 23'h00_0000;
  assign high_exp__380 = 8'hff;
  assign result_fraction__786 = 23'h00_0000;
  assign ne_171615 = x_fraction__142 != result_fraction__787;
  assign ne_171617 = prod_fraction__51 != result_fraction__788;
  assign eq_171618 = x_bexp__284 == high_exp__197;
  assign eq_171619 = x_fraction__284 == result_fraction__597;
  assign eq_171620 = prod_bexp__140 == high_exp__198;
  assign eq_171621 = prod_fraction__104 == result_fraction__598;
  assign high_exp__411 = 8'hff;
  assign result_fraction__818 = 23'h00_0000;
  assign high_exp__412 = 8'hff;
  assign result_fraction__819 = 23'h00_0000;
  assign ne_171633 = x_fraction__283 != result_fraction__820;
  assign ne_171635 = prod_fraction__103 != result_fraction__821;
  assign eq_171636 = x_bexp__428 == high_exp__265;
  assign eq_171637 = x_fraction__428 == result_fraction__664;
  assign eq_171638 = prod_bexp__212 == high_exp__266;
  assign eq_171639 = prod_fraction__158 == result_fraction__665;
  assign high_exp__443 = 8'hff;
  assign result_fraction__851 = 23'h00_0000;
  assign high_exp__444 = 8'hff;
  assign result_fraction__852 = 23'h00_0000;
  assign ne_171651 = x_fraction__427 != result_fraction__853;
  assign ne_171653 = prod_fraction__157 != result_fraction__854;
  assign eq_171654 = x_bexp__572 == high_exp__339;
  assign eq_171655 = x_fraction__572 == result_fraction__743;
  assign eq_171656 = prod_bexp__284 == high_exp__340;
  assign eq_171657 = prod_fraction__212 == result_fraction__744;
  assign high_exp__475 = 8'hff;
  assign result_fraction__884 = 23'h00_0000;
  assign high_exp__476 = 8'hff;
  assign result_fraction__885 = 23'h00_0000;
  assign ne_171669 = x_fraction__571 != result_fraction__886;
  assign ne_171671 = prod_fraction__211 != result_fraction__887;
  assign ne_171678 = x_fraction__70 != result_fraction__785;
  assign ne_171680 = prod_fraction__25 != result_fraction__786;
  assign fraction_shift__382 = 3'h3;
  assign fraction_shift__259 = 3'h4;
  assign is_operand_inf__17 = eq_171549 & eq_171550 | eq_171551 & eq_171552;
  assign and_reduce_171685 = &wide_exponent__53[7:0];
  assign ne_171697 = x_fraction__284 != result_fraction__818;
  assign ne_171699 = prod_fraction__104 != result_fraction__819;
  assign fraction_shift__400 = 3'h3;
  assign fraction_shift__294 = 3'h4;
  assign is_operand_inf__36 = eq_171563 & eq_171564 | eq_171565 & eq_171566;
  assign and_reduce_171704 = &wide_exponent__110[7:0];
  assign ne_171716 = x_fraction__428 != result_fraction__851;
  assign ne_171718 = prod_fraction__158 != result_fraction__852;
  assign fraction_shift__418 = 3'h3;
  assign fraction_shift__329 = 3'h4;
  assign is_operand_inf__55 = eq_171577 & eq_171578 | eq_171579 & eq_171580;
  assign and_reduce_171723 = &wide_exponent__167[7:0];
  assign ne_171735 = x_fraction__572 != result_fraction__884;
  assign ne_171737 = prod_fraction__212 != result_fraction__885;
  assign fraction_shift__436 = 3'h3;
  assign fraction_shift__364 = 3'h4;
  assign is_operand_inf__74 = eq_171591 & eq_171592 | eq_171593 & eq_171594;
  assign and_reduce_171742 = &wide_exponent__224[7:0];
  assign fraction_shift__383 = 3'h3;
  assign fraction_shift__260 = 3'h4;
  assign is_operand_inf__18 = eq_171600 & eq_171601 | eq_171602 & eq_171603;
  assign and_reduce_171752 = &wide_exponent__54[7:0];
  assign fraction_shift__54 = rounding_carry__17 ? fraction_shift__259 : fraction_shift__382;
  assign has_pos_inf__17 = ~(x_bexp__142 != high_exp__381 | ne_171615 | x_sign__36) | ~(prod_bexp__70 != high_exp__382 | ne_171617 | prod_sign__17);
  assign has_neg_inf__17 = eq_171549 & eq_171550 & x_sign__36 | eq_171551 & eq_171552 & prod_sign__17;
  assign fraction_shift__401 = 3'h3;
  assign fraction_shift__295 = 3'h4;
  assign is_operand_inf__37 = eq_171618 & eq_171619 | eq_171620 & eq_171621;
  assign and_reduce_171766 = &wide_exponent__111[7:0];
  assign fraction_shift__110 = rounding_carry__36 ? fraction_shift__294 : fraction_shift__400;
  assign has_pos_inf__36 = ~(x_bexp__283 != high_exp__413 | ne_171633 | x_sign__71) | ~(prod_bexp__139 != high_exp__414 | ne_171635 | prod_sign__35);
  assign has_neg_inf__36 = eq_171563 & eq_171564 & x_sign__71 | eq_171565 & eq_171566 & prod_sign__35;
  assign fraction_shift__419 = 3'h3;
  assign fraction_shift__330 = 3'h4;
  assign is_operand_inf__56 = eq_171636 & eq_171637 | eq_171638 & eq_171639;
  assign and_reduce_171780 = &wide_exponent__168[7:0];
  assign fraction_shift__167 = rounding_carry__55 ? fraction_shift__329 : fraction_shift__418;
  assign has_pos_inf__55 = ~(x_bexp__427 != high_exp__445 | ne_171651 | x_sign__107) | ~(prod_bexp__211 != high_exp__446 | ne_171653 | prod_sign__53);
  assign has_neg_inf__55 = eq_171577 & eq_171578 & x_sign__107 | eq_171579 & eq_171580 & prod_sign__53;
  assign fraction_shift__437 = 3'h3;
  assign fraction_shift__365 = 3'h4;
  assign is_operand_inf__75 = eq_171654 & eq_171655 | eq_171656 & eq_171657;
  assign and_reduce_171794 = &wide_exponent__225[7:0];
  assign fraction_shift__224 = rounding_carry__74 ? fraction_shift__364 : fraction_shift__436;
  assign has_pos_inf__74 = ~(x_bexp__571 != high_exp__477 | ne_171669 | x_sign__143) | ~(prod_bexp__283 != high_exp__478 | ne_171671 | prod_sign__71);
  assign has_neg_inf__74 = eq_171591 & eq_171592 & x_sign__143 | eq_171593 & eq_171594 & prod_sign__71;
  assign fraction_shift__27 = rounding_carry__18 ? fraction_shift__260 : fraction_shift__383;
  assign has_pos_inf__18 = ~(x_bexp__70 != high_exp__379 | ne_171678 | x_sign__18) | ~(prod_bexp__34 != high_exp__380 | ne_171680 | prod_sign__18);
  assign has_neg_inf__18 = eq_171600 & eq_171601 & x_sign__18 | eq_171602 & eq_171603 & prod_sign__18;
  assign shrl_171808 = rounded_fraction__17 >> fraction_shift__54;
  assign fraction_shift__111 = rounding_carry__37 ? fraction_shift__295 : fraction_shift__401;
  assign has_pos_inf__37 = ~(x_bexp__284 != high_exp__411 | ne_171697 | x_sign__72) | ~(prod_bexp__140 != high_exp__412 | ne_171699 | prod_sign__36);
  assign has_neg_inf__37 = eq_171618 & eq_171619 & x_sign__72 | eq_171620 & eq_171621 & prod_sign__36;
  assign shrl_171817 = rounded_fraction__36 >> fraction_shift__110;
  assign fraction_shift__168 = rounding_carry__56 ? fraction_shift__330 : fraction_shift__419;
  assign has_pos_inf__56 = ~(x_bexp__428 != high_exp__443 | ne_171716 | x_sign__108) | ~(prod_bexp__212 != high_exp__444 | ne_171718 | prod_sign__54);
  assign has_neg_inf__56 = eq_171636 & eq_171637 & x_sign__108 | eq_171638 & eq_171639 & prod_sign__54;
  assign shrl_171826 = rounded_fraction__55 >> fraction_shift__167;
  assign fraction_shift__225 = rounding_carry__75 ? fraction_shift__365 : fraction_shift__437;
  assign has_pos_inf__75 = ~(x_bexp__572 != high_exp__475 | ne_171735 | x_sign__144) | ~(prod_bexp__284 != high_exp__476 | ne_171737 | prod_sign__72);
  assign has_neg_inf__75 = eq_171654 & eq_171655 & x_sign__144 | eq_171656 & eq_171657 & prod_sign__72;
  assign shrl_171835 = rounded_fraction__74 >> fraction_shift__224;
  assign shrl_171840 = rounded_fraction__18 >> fraction_shift__27;
  assign result_fraction__105 = shrl_171808[22:0];
  assign is_result_nan__35 = eq_171549 & ne_171615 | eq_171551 & ne_171617 | has_pos_inf__17 & has_neg_inf__17;
  assign shrl_171848 = rounded_fraction__37 >> fraction_shift__111;
  assign result_fraction__220 = shrl_171817[22:0];
  assign is_result_nan__74 = eq_171563 & ne_171633 | eq_171565 & ne_171635 | has_pos_inf__36 & has_neg_inf__36;
  assign shrl_171856 = rounded_fraction__56 >> fraction_shift__168;
  assign result_fraction__337 = shrl_171826[22:0];
  assign is_result_nan__113 = eq_171577 & ne_171651 | eq_171579 & ne_171653 | has_pos_inf__55 & has_neg_inf__55;
  assign shrl_171864 = rounded_fraction__75 >> fraction_shift__225;
  assign result_fraction__454 = shrl_171835[22:0];
  assign is_result_nan__152 = eq_171591 & ne_171669 | eq_171593 & ne_171671 | has_pos_inf__74 & has_neg_inf__74;
  assign result_fraction__52 = shrl_171840[22:0];
  assign is_result_nan__36 = eq_171600 & ne_171678 | eq_171602 & ne_171680 | has_pos_inf__18 & has_neg_inf__18;
  assign result_fraction__106 = result_fraction__105 & {23{~(is_operand_inf__17 | wide_exponent__53[8] | and_reduce_171685 | ~((|wide_exponent__53[8:1]) | wide_exponent__53[0]))}};
  assign nan_fraction__101 = 23'h40_0000;
  assign or_171877 = is_result_nan__35 | is_operand_inf__17 | wide_exponent__53[8] | and_reduce_171685;
  assign high_exp__134 = 8'hff;
  assign result_fraction__221 = shrl_171848[22:0];
  assign is_result_nan__75 = eq_171618 & ne_171697 | eq_171620 & ne_171699 | has_pos_inf__37 & has_neg_inf__37;
  assign result_fraction__222 = result_fraction__220 & {23{~(is_operand_inf__36 | wide_exponent__110[8] | and_reduce_171704 | ~((|wide_exponent__110[8:1]) | wide_exponent__110[0]))}};
  assign nan_fraction__128 = 23'h40_0000;
  assign high_exp__199 = 8'hff;
  assign result_fraction__338 = shrl_171856[22:0];
  assign is_result_nan__114 = eq_171636 & ne_171716 | eq_171638 & ne_171718 | has_pos_inf__56 & has_neg_inf__56;
  assign result_fraction__339 = result_fraction__337 & {23{~(is_operand_inf__55 | wide_exponent__167[8] | and_reduce_171723 | ~((|wide_exponent__167[8:1]) | wide_exponent__167[0]))}};
  assign nan_fraction__157 = 23'h40_0000;
  assign high_exp__267 = 8'hff;
  assign result_fraction__455 = shrl_171864[22:0];
  assign is_result_nan__153 = eq_171654 & ne_171735 | eq_171656 & ne_171737 | has_pos_inf__75 & has_neg_inf__75;
  assign result_fraction__456 = result_fraction__454 & {23{~(is_operand_inf__74 | wide_exponent__224[8] | and_reduce_171742 | ~((|wide_exponent__224[8:1]) | wide_exponent__224[0]))}};
  assign nan_fraction__186 = 23'h40_0000;
  assign high_exp__341 = 8'hff;
  assign result_fraction__53 = result_fraction__52 & {23{~(is_operand_inf__18 | wide_exponent__54[8] | and_reduce_171752 | ~((|wide_exponent__54[8:1]) | wide_exponent__54[0]))}};
  assign nan_fraction__102 = 23'h40_0000;
  assign or_171902 = is_result_nan__36 | is_operand_inf__18 | wide_exponent__54[8] | and_reduce_171752;
  assign high_exp__135 = 8'hff;
  assign result_sign__466 = 1'h0;
  assign result_fraction__107 = is_result_nan__35 ? nan_fraction__101 : result_fraction__106;
  assign result_exponent__18 = or_171877 ? high_exp__134 : wide_exponent__53[7:0];
  assign x_bexp__812 = 8'h00;
  assign result_fraction__223 = result_fraction__221 & {23{~(is_operand_inf__37 | wide_exponent__111[8] | and_reduce_171766 | ~((|wide_exponent__111[8:1]) | wide_exponent__111[0]))}};
  assign nan_fraction__129 = 23'h40_0000;
  assign or_171910 = is_result_nan__75 | is_operand_inf__37 | wide_exponent__111[8] | and_reduce_171766;
  assign high_exp__200 = 8'hff;
  assign result_sign__563 = 1'h0;
  assign result_fraction__224 = is_result_nan__74 ? nan_fraction__128 : result_fraction__222;
  assign result_exponent__36 = is_result_nan__74 | is_operand_inf__36 | wide_exponent__110[8] | and_reduce_171704 ? high_exp__199 : wide_exponent__110[7:0];
  assign x_bexp__813 = 8'h00;
  assign result_fraction__340 = result_fraction__338 & {23{~(is_operand_inf__56 | wide_exponent__168[8] | and_reduce_171780 | ~((|wide_exponent__168[8:1]) | wide_exponent__168[0]))}};
  assign nan_fraction__158 = 23'h40_0000;
  assign or_171918 = is_result_nan__114 | is_operand_inf__56 | wide_exponent__168[8] | and_reduce_171780;
  assign high_exp__268 = 8'hff;
  assign result_sign__665 = 1'h0;
  assign result_fraction__341 = is_result_nan__113 ? nan_fraction__157 : result_fraction__339;
  assign result_exponent__55 = is_result_nan__113 | is_operand_inf__55 | wide_exponent__167[8] | and_reduce_171723 ? high_exp__267 : wide_exponent__167[7:0];
  assign x_bexp__814 = 8'h00;
  assign result_fraction__457 = result_fraction__455 & {23{~(is_operand_inf__75 | wide_exponent__225[8] | and_reduce_171794 | ~((|wide_exponent__225[8:1]) | wide_exponent__225[0]))}};
  assign nan_fraction__187 = 23'h40_0000;
  assign or_171926 = is_result_nan__153 | is_operand_inf__75 | wide_exponent__225[8] | and_reduce_171794;
  assign high_exp__342 = 8'hff;
  assign result_sign__777 = 1'h0;
  assign result_fraction__458 = is_result_nan__152 ? nan_fraction__186 : result_fraction__456;
  assign result_exponent__74 = is_result_nan__152 | is_operand_inf__74 | wide_exponent__224[8] | and_reduce_171742 ? high_exp__341 : wide_exponent__224[7:0];
  assign x_bexp__815 = 8'h00;
  assign result_sign__467 = 1'h0;
  assign result_fraction__108 = is_result_nan__36 ? nan_fraction__102 : result_fraction__53;
  assign result_exponent__9 = or_171902 ? high_exp__135 : wide_exponent__54[7:0];
  assign x_bexp__816 = 8'h00;
  assign ne_171938 = result_exponent__18 != x_bexp__812;
  assign result_sign__564 = 1'h0;
  assign result_fraction__225 = is_result_nan__75 ? nan_fraction__129 : result_fraction__223;
  assign result_exponent__37 = or_171910 ? high_exp__200 : wide_exponent__111[7:0];
  assign x_bexp__817 = 8'h00;
  assign ne_171945 = result_exponent__36 != x_bexp__813;
  assign result_sign__666 = 1'h0;
  assign result_fraction__342 = is_result_nan__114 ? nan_fraction__158 : result_fraction__340;
  assign result_exponent__56 = or_171918 ? high_exp__268 : wide_exponent__168[7:0];
  assign x_bexp__818 = 8'h00;
  assign ne_171952 = result_exponent__55 != x_bexp__814;
  assign result_sign__778 = 1'h0;
  assign result_fraction__459 = is_result_nan__153 ? nan_fraction__187 : result_fraction__457;
  assign result_exponent__75 = or_171926 ? high_exp__342 : wide_exponent__225[7:0];
  assign x_bexp__819 = 8'h00;
  assign ne_171959 = result_exponent__74 != x_bexp__815;
  assign ne_171962 = result_exponent__9 != x_bexp__816;
  assign result_sign__468 = 1'h0;
  assign y_stencil_out_fraction__5 = {result_sign__466, result_fraction__107} | 24'h80_0000;
  assign ne_171968 = result_exponent__37 != x_bexp__817;
  assign result_sign__565 = 1'h0;
  assign y_stencil_out_fraction__13 = {result_sign__563, result_fraction__224} | 24'h80_0000;
  assign ne_171974 = result_exponent__56 != x_bexp__818;
  assign result_sign__667 = 1'h0;
  assign y_stencil_out_fraction__23 = {result_sign__665, result_fraction__341} | 24'h80_0000;
  assign ne_171980 = result_exponent__75 != x_bexp__819;
  assign result_sign__779 = 1'h0;
  assign y_stencil_out_fraction__33 = {result_sign__777, result_fraction__458} | 24'h80_0000;
  assign result_sign__469 = 1'h0;
  assign x_stencil_out_fraction__5 = {result_sign__467, result_fraction__108} | 24'h80_0000;
  assign y_stencil_out_fraction__3 = y_stencil_out_fraction__5 & {24{ne_171938}};
  assign result_sign__566 = 1'h0;
  assign x_stencil_out_fraction__13 = {result_sign__564, result_fraction__225} | 24'h80_0000;
  assign y_stencil_out_fraction__15 = y_stencil_out_fraction__13 & {24{ne_171945}};
  assign result_sign__668 = 1'h0;
  assign x_stencil_out_fraction__23 = {result_sign__666, result_fraction__342} | 24'h80_0000;
  assign y_stencil_out_fraction__25 = y_stencil_out_fraction__23 & {24{ne_171952}};
  assign result_sign__780 = 1'h0;
  assign x_stencil_out_fraction__33 = {result_sign__778, result_fraction__459} | 24'h80_0000;
  assign y_stencil_out_fraction__35 = y_stencil_out_fraction__33 & {24{ne_171959}};
  assign x_stencil_out_fraction__3 = x_stencil_out_fraction__5 & {24{ne_171962}};
  assign result_sign__470 = 1'h0;
  assign add_172007 = {result_sign__468, result_exponent__18} + {result_sign__468, result_exponent__18};
  assign fraction__170 = umul48b_24b_x_24b(y_stencil_out_fraction__3, y_stencil_out_fraction__3);
  assign x_stencil_out_fraction__15 = x_stencil_out_fraction__13 & {24{ne_171968}};
  assign result_sign__567 = 1'h0;
  assign add_172012 = {result_sign__565, result_exponent__36} + {result_sign__565, result_exponent__36};
  assign fraction__342 = umul48b_24b_x_24b(y_stencil_out_fraction__15, y_stencil_out_fraction__15);
  assign x_stencil_out_fraction__25 = x_stencil_out_fraction__23 & {24{ne_171974}};
  assign result_sign__669 = 1'h0;
  assign add_172017 = {result_sign__667, result_exponent__55} + {result_sign__667, result_exponent__55};
  assign fraction__521 = umul48b_24b_x_24b(y_stencil_out_fraction__25, y_stencil_out_fraction__25);
  assign x_stencil_out_fraction__35 = x_stencil_out_fraction__33 & {24{ne_171980}};
  assign result_sign__781 = 1'h0;
  assign add_172022 = {result_sign__779, result_exponent__74} + {result_sign__779, result_exponent__74};
  assign fraction__700 = umul48b_24b_x_24b(y_stencil_out_fraction__35, y_stencil_out_fraction__35);
  assign result_sign__471 = 1'h0;
  assign add_172025 = {result_sign__469, result_exponent__9} + {result_sign__469, result_exponent__9};
  assign fraction__163 = umul48b_24b_x_24b(x_stencil_out_fraction__3, x_stencil_out_fraction__3);
  assign result_sign__568 = 1'h0;
  assign add_172033 = {result_sign__566, result_exponent__37} + {result_sign__566, result_exponent__37};
  assign fraction__343 = umul48b_24b_x_24b(x_stencil_out_fraction__15, x_stencil_out_fraction__15);
  assign result_sign__670 = 1'h0;
  assign add_172041 = {result_sign__668, result_exponent__56} + {result_sign__668, result_exponent__56};
  assign fraction__522 = umul48b_24b_x_24b(x_stencil_out_fraction__25, x_stencil_out_fraction__25);
  assign result_sign__782 = 1'h0;
  assign add_172049 = {result_sign__780, result_exponent__75} + {result_sign__780, result_exponent__75};
  assign fraction__701 = umul48b_24b_x_24b(x_stencil_out_fraction__35, x_stencil_out_fraction__35);
  assign exp__76 = {result_sign__470, add_172007} + 10'h381;
  assign fraction__171 = fraction__170 >> fraction__170[47];
  assign sticky__56 = {47'h0000_0000_0000, fraction__170[0]};
  assign exp__155 = {result_sign__567, add_172012} + 10'h381;
  assign fraction__344 = fraction__342 >> fraction__342[47];
  assign sticky__114 = {47'h0000_0000_0000, fraction__342[0]};
  assign exp__237 = {result_sign__669, add_172017} + 10'h381;
  assign fraction__523 = fraction__521 >> fraction__521[47];
  assign sticky__173 = {47'h0000_0000_0000, fraction__521[0]};
  assign exp__319 = {result_sign__781, add_172022} + 10'h381;
  assign fraction__702 = fraction__700 >> fraction__700[47];
  assign sticky__232 = {47'h0000_0000_0000, fraction__700[0]};
  assign exp__73 = {result_sign__471, add_172025} + 10'h381;
  assign fraction__164 = fraction__163 >> fraction__163[47];
  assign sticky__55 = {47'h0000_0000_0000, fraction__163[0]};
  assign exp__77 = exp__76 & {10{ne_171938}};
  assign fraction__172 = fraction__171 | sticky__56;
  assign exp__156 = {result_sign__568, add_172033} + 10'h381;
  assign fraction__345 = fraction__343 >> fraction__343[47];
  assign sticky__115 = {47'h0000_0000_0000, fraction__343[0]};
  assign exp__157 = exp__155 & {10{ne_171945}};
  assign fraction__346 = fraction__344 | sticky__114;
  assign exp__238 = {result_sign__670, add_172041} + 10'h381;
  assign fraction__524 = fraction__522 >> fraction__522[47];
  assign sticky__174 = {47'h0000_0000_0000, fraction__522[0]};
  assign exp__239 = exp__237 & {10{ne_171952}};
  assign fraction__525 = fraction__523 | sticky__173;
  assign exp__320 = {result_sign__782, add_172049} + 10'h381;
  assign fraction__703 = fraction__701 >> fraction__701[47];
  assign sticky__233 = {47'h0000_0000_0000, fraction__701[0]};
  assign exp__321 = exp__319 & {10{ne_171959}};
  assign fraction__704 = fraction__702 | sticky__232;
  assign exp__74 = exp__73 & {10{ne_171962}};
  assign fraction__165 = fraction__164 | sticky__55;
  assign exp__78 = exp__77 + {9'h000, fraction__170[47]};
  assign result_sign__472 = 1'h0;
  assign exp__158 = exp__156 & {10{ne_171968}};
  assign fraction__347 = fraction__345 | sticky__115;
  assign exp__159 = exp__157 + {9'h000, fraction__342[47]};
  assign result_sign__569 = 1'h0;
  assign exp__240 = exp__238 & {10{ne_171974}};
  assign fraction__526 = fraction__524 | sticky__174;
  assign exp__241 = exp__239 + {9'h000, fraction__521[47]};
  assign result_sign__671 = 1'h0;
  assign exp__322 = exp__320 & {10{ne_171980}};
  assign fraction__705 = fraction__703 | sticky__233;
  assign exp__323 = exp__321 + {9'h000, fraction__700[47]};
  assign result_sign__783 = 1'h0;
  assign exp__75 = exp__74 + {9'h000, fraction__163[47]};
  assign result_sign__473 = 1'h0;
  assign exp__160 = exp__158 + {9'h000, fraction__343[47]};
  assign result_sign__570 = 1'h0;
  assign exp__242 = exp__240 + {9'h000, fraction__522[47]};
  assign result_sign__672 = 1'h0;
  assign exp__324 = exp__322 + {9'h000, fraction__701[47]};
  assign result_sign__784 = 1'h0;
  assign fraction__173 = $signed(exp__78) <= $signed(10'h000) ? {result_sign__472, fraction__172[47:1]} : fraction__172;
  assign sticky__57 = {47'h0000_0000_0000, fraction__172[0]};
  assign fraction__348 = $signed(exp__159) <= $signed(10'h000) ? {result_sign__569, fraction__346[47:1]} : fraction__346;
  assign sticky__116 = {47'h0000_0000_0000, fraction__346[0]};
  assign fraction__527 = $signed(exp__241) <= $signed(10'h000) ? {result_sign__671, fraction__525[47:1]} : fraction__525;
  assign sticky__175 = {47'h0000_0000_0000, fraction__525[0]};
  assign fraction__706 = $signed(exp__323) <= $signed(10'h000) ? {result_sign__783, fraction__704[47:1]} : fraction__704;
  assign sticky__234 = {47'h0000_0000_0000, fraction__704[0]};
  assign fraction__166 = $signed(exp__75) <= $signed(10'h000) ? {result_sign__473, fraction__165[47:1]} : fraction__165;
  assign sticky__58 = {47'h0000_0000_0000, fraction__165[0]};
  assign fraction__174 = fraction__173 | sticky__57;
  assign fraction__349 = $signed(exp__160) <= $signed(10'h000) ? {result_sign__570, fraction__347[47:1]} : fraction__347;
  assign sticky__117 = {47'h0000_0000_0000, fraction__347[0]};
  assign fraction__350 = fraction__348 | sticky__116;
  assign fraction__528 = $signed(exp__242) <= $signed(10'h000) ? {result_sign__672, fraction__526[47:1]} : fraction__526;
  assign sticky__176 = {47'h0000_0000_0000, fraction__526[0]};
  assign fraction__529 = fraction__527 | sticky__175;
  assign fraction__707 = $signed(exp__324) <= $signed(10'h000) ? {result_sign__784, fraction__705[47:1]} : fraction__705;
  assign sticky__235 = {47'h0000_0000_0000, fraction__705[0]};
  assign fraction__708 = fraction__706 | sticky__234;
  assign fraction__167 = fraction__166 | sticky__58;
  assign fraction__351 = fraction__349 | sticky__117;
  assign fraction__530 = fraction__528 | sticky__176;
  assign fraction__709 = fraction__707 | sticky__235;
  assign result_sign__474 = 1'h0;
  assign fraction__175 = fraction__174[45:23];
  assign result_sign__571 = 1'h0;
  assign fraction__352 = fraction__350[45:23];
  assign result_sign__673 = 1'h0;
  assign fraction__531 = fraction__529[45:23];
  assign result_sign__785 = 1'h0;
  assign fraction__710 = fraction__708[45:23];
  assign result_sign__475 = 1'h0;
  assign fraction__168 = fraction__167[45:23];
  assign greater_than_half_way__19 = fraction__174[22] & fraction__174[21:0] != 22'h00_0000;
  assign fraction__176 = {result_sign__474, fraction__175};
  assign result_sign__572 = 1'h0;
  assign fraction__353 = fraction__351[45:23];
  assign greater_than_half_way__39 = fraction__350[22] & fraction__350[21:0] != 22'h00_0000;
  assign fraction__354 = {result_sign__571, fraction__352};
  assign result_sign__674 = 1'h0;
  assign fraction__532 = fraction__530[45:23];
  assign greater_than_half_way__59 = fraction__529[22] & fraction__529[21:0] != 22'h00_0000;
  assign fraction__533 = {result_sign__673, fraction__531};
  assign result_sign__786 = 1'h0;
  assign fraction__711 = fraction__709[45:23];
  assign greater_than_half_way__79 = fraction__708[22] & fraction__708[21:0] != 22'h00_0000;
  assign fraction__712 = {result_sign__785, fraction__710};
  assign greater_than_half_way__20 = fraction__167[22] & fraction__167[21:0] != 22'h00_0000;
  assign fraction__169 = {result_sign__475, fraction__168};
  assign do_round_up__37 = greater_than_half_way__19 | fraction__174[22] & fraction__174[21:0] == 22'h00_0000 & fraction__174[23];
  assign add_172321 = fraction__176 + 24'h00_0001;
  assign greater_than_half_way__40 = fraction__351[22] & fraction__351[21:0] != 22'h00_0000;
  assign fraction__355 = {result_sign__572, fraction__353};
  assign do_round_up__76 = greater_than_half_way__39 | fraction__350[22] & fraction__350[21:0] == 22'h00_0000 & fraction__350[23];
  assign add_172327 = fraction__354 + 24'h00_0001;
  assign greater_than_half_way__60 = fraction__530[22] & fraction__530[21:0] != 22'h00_0000;
  assign fraction__534 = {result_sign__674, fraction__532};
  assign do_round_up__115 = greater_than_half_way__59 | fraction__529[22] & fraction__529[21:0] == 22'h00_0000 & fraction__529[23];
  assign add_172333 = fraction__533 + 24'h00_0001;
  assign greater_than_half_way__80 = fraction__709[22] & fraction__709[21:0] != 22'h00_0000;
  assign fraction__713 = {result_sign__786, fraction__711};
  assign do_round_up__154 = greater_than_half_way__79 | fraction__708[22] & fraction__708[21:0] == 22'h00_0000 & fraction__708[23];
  assign add_172339 = fraction__712 + 24'h00_0001;
  assign do_round_up__38 = greater_than_half_way__20 | fraction__167[22] & fraction__167[21:0] == 22'h00_0000 & fraction__167[23];
  assign add_172341 = fraction__169 + 24'h00_0001;
  assign fraction__177 = do_round_up__37 ? add_172321 : fraction__176;
  assign do_round_up__77 = greater_than_half_way__40 | fraction__351[22] & fraction__351[21:0] == 22'h00_0000 & fraction__351[23];
  assign add_172345 = fraction__355 + 24'h00_0001;
  assign fraction__356 = do_round_up__76 ? add_172327 : fraction__354;
  assign do_round_up__116 = greater_than_half_way__60 | fraction__530[22] & fraction__530[21:0] == 22'h00_0000 & fraction__530[23];
  assign add_172349 = fraction__534 + 24'h00_0001;
  assign fraction__535 = do_round_up__115 ? add_172333 : fraction__533;
  assign do_round_up__155 = greater_than_half_way__80 | fraction__709[22] & fraction__709[21:0] == 22'h00_0000 & fraction__709[23];
  assign add_172353 = fraction__713 + 24'h00_0001;
  assign fraction__714 = do_round_up__154 ? add_172339 : fraction__712;
  assign fraction__178 = do_round_up__38 ? add_172341 : fraction__169;
  assign add_172359 = exp__78 + 10'h001;
  assign fraction__357 = do_round_up__77 ? add_172345 : fraction__355;
  assign add_172363 = exp__159 + 10'h001;
  assign fraction__536 = do_round_up__116 ? add_172349 : fraction__534;
  assign add_172367 = exp__241 + 10'h001;
  assign fraction__715 = do_round_up__155 ? add_172353 : fraction__713;
  assign add_172371 = exp__323 + 10'h001;
  assign add_172373 = exp__75 + 10'h001;
  assign exp__79 = fraction__177[23] ? add_172359 : exp__78;
  assign add_172377 = exp__160 + 10'h001;
  assign exp__161 = fraction__356[23] ? add_172363 : exp__159;
  assign add_172381 = exp__242 + 10'h001;
  assign exp__243 = fraction__535[23] ? add_172367 : exp__241;
  assign add_172385 = exp__324 + 10'h001;
  assign exp__325 = fraction__714[23] ? add_172371 : exp__323;
  assign exp__80 = fraction__178[23] ? add_172373 : exp__75;
  assign exp__162 = fraction__357[23] ? add_172377 : exp__160;
  assign exp__244 = fraction__536[23] ? add_172381 : exp__242;
  assign exp__326 = fraction__715[23] ? add_172385 : exp__324;
  assign result_exp__57 = exp__79[8:0];
  assign result_exp__115 = exp__161[8:0];
  assign result_exp__175 = exp__243[8:0];
  assign result_exp__235 = exp__325[8:0];
  assign result_exp__55 = exp__80[8:0];
  assign result_fraction__534 = 23'h00_0000;
  assign result_fraction__532 = 23'h00_0000;
  assign result_exp__58 = result_exp__57 & {9{$signed(exp__79) > $signed(10'h000)}};
  assign result_exp__116 = exp__162[8:0];
  assign high_exp__201 = 8'hff;
  assign result_fraction__601 = 23'h00_0000;
  assign result_fraction__599 = 23'h00_0000;
  assign result_exp__117 = result_exp__115 & {9{$signed(exp__161) > $signed(10'h000)}};
  assign result_exp__176 = exp__244[8:0];
  assign high_exp__269 = 8'hff;
  assign result_fraction__668 = 23'h00_0000;
  assign result_fraction__666 = 23'h00_0000;
  assign result_exp__177 = result_exp__175 & {9{$signed(exp__243) > $signed(10'h000)}};
  assign result_exp__236 = exp__326[8:0];
  assign high_exp__343 = 8'hff;
  assign result_fraction__747 = 23'h00_0000;
  assign result_fraction__745 = 23'h00_0000;
  assign result_exp__237 = result_exp__235 & {9{$signed(exp__325) > $signed(10'h000)}};
  assign result_fraction__535 = 23'h00_0000;
  assign result_fraction__533 = 23'h00_0000;
  assign result_exp__56 = result_exp__55 & {9{$signed(exp__80) > $signed(10'h000)}};
  assign result_fraction__602 = 23'h00_0000;
  assign result_fraction__600 = 23'h00_0000;
  assign result_exp__118 = result_exp__116 & {9{$signed(exp__162) > $signed(10'h000)}};
  assign eq_172444 = result_exponent__36 == high_exp__201;
  assign result_fraction__669 = 23'h00_0000;
  assign result_fraction__667 = 23'h00_0000;
  assign result_exp__178 = result_exp__176 & {9{$signed(exp__244) > $signed(10'h000)}};
  assign eq_172451 = result_exponent__55 == high_exp__269;
  assign result_fraction__748 = 23'h00_0000;
  assign result_fraction__746 = 23'h00_0000;
  assign result_exp__238 = result_exp__236 & {9{$signed(exp__326) > $signed(10'h000)}};
  assign eq_172458 = result_exponent__74 == high_exp__343;
  assign is_result_nan__37 = or_171877 & result_fraction__107 != result_fraction__534;
  assign has_inf_arg__19 = or_171877 & result_fraction__107 == result_fraction__532;
  assign and_reduce_172468 = &result_exp__58[7:0];
  assign is_result_nan__76 = eq_172444 & result_fraction__224 != result_fraction__601;
  assign has_inf_arg__39 = eq_172444 & result_fraction__224 == result_fraction__599;
  assign and_reduce_172475 = &result_exp__117[7:0];
  assign is_result_nan__115 = eq_172451 & result_fraction__341 != result_fraction__668;
  assign has_inf_arg__59 = eq_172451 & result_fraction__341 == result_fraction__666;
  assign and_reduce_172482 = &result_exp__177[7:0];
  assign is_result_nan__154 = eq_172458 & result_fraction__458 != result_fraction__747;
  assign has_inf_arg__79 = eq_172458 & result_fraction__458 == result_fraction__745;
  assign and_reduce_172489 = &result_exp__237[7:0];
  assign is_result_nan__38 = or_171902 & result_fraction__108 != result_fraction__535;
  assign has_inf_arg__20 = or_171902 & result_fraction__108 == result_fraction__533;
  assign and_reduce_172495 = &result_exp__56[7:0];
  assign high_exp__136 = 8'hff;
  assign is_result_nan__77 = or_171910 & result_fraction__225 != result_fraction__602;
  assign has_inf_arg__40 = or_171910 & result_fraction__225 == result_fraction__600;
  assign and_reduce_172503 = &result_exp__118[7:0];
  assign high_exp__202 = 8'hff;
  assign is_result_nan__116 = or_171918 & result_fraction__342 != result_fraction__669;
  assign has_inf_arg__60 = or_171918 & result_fraction__342 == result_fraction__667;
  assign and_reduce_172511 = &result_exp__178[7:0];
  assign high_exp__270 = 8'hff;
  assign is_result_nan__155 = or_171926 & result_fraction__459 != result_fraction__748;
  assign has_inf_arg__80 = or_171926 & result_fraction__459 == result_fraction__746;
  assign and_reduce_172519 = &result_exp__238[7:0];
  assign high_exp__344 = 8'hff;
  assign is_subnormal__20 = $signed(exp__80) <= $signed(10'h000);
  assign is_subnormal__19 = $signed(exp__79) <= $signed(10'h000);
  assign high_exp__137 = 8'hff;
  assign result_exp__59 = is_result_nan__37 | has_inf_arg__19 | result_exp__58[8] | and_reduce_172468 ? high_exp__136 : result_exp__58[7:0];
  assign is_subnormal__40 = $signed(exp__162) <= $signed(10'h000);
  assign is_subnormal__39 = $signed(exp__161) <= $signed(10'h000);
  assign high_exp__203 = 8'hff;
  assign result_exp__119 = is_result_nan__76 | has_inf_arg__39 | result_exp__117[8] | and_reduce_172475 ? high_exp__202 : result_exp__117[7:0];
  assign is_subnormal__60 = $signed(exp__244) <= $signed(10'h000);
  assign is_subnormal__59 = $signed(exp__243) <= $signed(10'h000);
  assign high_exp__271 = 8'hff;
  assign result_exp__179 = is_result_nan__115 | has_inf_arg__59 | result_exp__177[8] | and_reduce_172482 ? high_exp__270 : result_exp__177[7:0];
  assign is_subnormal__80 = $signed(exp__326) <= $signed(10'h000);
  assign is_subnormal__79 = $signed(exp__325) <= $signed(10'h000);
  assign high_exp__345 = 8'hff;
  assign result_exp__239 = is_result_nan__154 | has_inf_arg__79 | result_exp__237[8] | and_reduce_172489 ? high_exp__344 : result_exp__237[7:0];
  assign result_sign__476 = 1'h0;
  assign result_exp__60 = is_result_nan__38 | has_inf_arg__20 | result_exp__56[8] | and_reduce_172495 ? high_exp__137 : result_exp__56[7:0];
  assign result_sign__477 = 1'h0;
  assign result_sign__573 = 1'h0;
  assign result_exp__120 = is_result_nan__77 | has_inf_arg__40 | result_exp__118[8] | and_reduce_172503 ? high_exp__203 : result_exp__118[7:0];
  assign result_sign__574 = 1'h0;
  assign result_sign__675 = 1'h0;
  assign result_exp__180 = is_result_nan__116 | has_inf_arg__60 | result_exp__178[8] | and_reduce_172511 ? high_exp__271 : result_exp__178[7:0];
  assign result_sign__676 = 1'h0;
  assign result_sign__787 = 1'h0;
  assign result_exp__240 = is_result_nan__155 | has_inf_arg__80 | result_exp__238[8] | and_reduce_172519 ? high_exp__345 : result_exp__238[7:0];
  assign result_sign__788 = 1'h0;
  assign result_fraction__109 = fraction__178[22:0];
  assign result_fraction__111 = fraction__177[22:0];
  assign sum__19 = {result_sign__476, result_exp__60} + {result_sign__477, ~result_exp__59};
  assign result_fraction__227 = fraction__357[22:0];
  assign result_fraction__226 = fraction__356[22:0];
  assign sum__38 = {result_sign__573, result_exp__120} + {result_sign__574, ~result_exp__119};
  assign result_fraction__344 = fraction__536[22:0];
  assign result_fraction__343 = fraction__535[22:0];
  assign sum__57 = {result_sign__675, result_exp__180} + {result_sign__676, ~result_exp__179};
  assign result_fraction__461 = fraction__715[22:0];
  assign result_fraction__460 = fraction__714[22:0];
  assign sum__76 = {result_sign__787, result_exp__240} + {result_sign__788, ~result_exp__239};
  assign result_fraction__110 = result_fraction__109 & {23{~(has_inf_arg__20 | result_exp__56[8] | and_reduce_172495 | is_subnormal__20)}};
  assign nan_fraction__104 = 23'h40_0000;
  assign result_fraction__112 = result_fraction__111 & {23{~(has_inf_arg__19 | result_exp__58[8] | and_reduce_172468 | is_subnormal__19)}};
  assign nan_fraction__103 = 23'h40_0000;
  assign result_fraction__229 = result_fraction__227 & {23{~(has_inf_arg__40 | result_exp__118[8] | and_reduce_172503 | is_subnormal__40)}};
  assign nan_fraction__131 = 23'h40_0000;
  assign result_fraction__228 = result_fraction__226 & {23{~(has_inf_arg__39 | result_exp__117[8] | and_reduce_172475 | is_subnormal__39)}};
  assign nan_fraction__130 = 23'h40_0000;
  assign result_fraction__346 = result_fraction__344 & {23{~(has_inf_arg__60 | result_exp__178[8] | and_reduce_172511 | is_subnormal__60)}};
  assign nan_fraction__160 = 23'h40_0000;
  assign result_fraction__345 = result_fraction__343 & {23{~(has_inf_arg__59 | result_exp__177[8] | and_reduce_172482 | is_subnormal__59)}};
  assign nan_fraction__159 = 23'h40_0000;
  assign result_fraction__463 = result_fraction__461 & {23{~(has_inf_arg__80 | result_exp__238[8] | and_reduce_172519 | is_subnormal__80)}};
  assign nan_fraction__189 = 23'h40_0000;
  assign result_fraction__462 = result_fraction__460 & {23{~(has_inf_arg__79 | result_exp__237[8] | and_reduce_172489 | is_subnormal__79)}};
  assign nan_fraction__188 = 23'h40_0000;
  assign result_fraction__114 = is_result_nan__38 ? nan_fraction__104 : result_fraction__110;
  assign result_fraction__113 = is_result_nan__37 ? nan_fraction__103 : result_fraction__112;
  assign y_sq_bexp__1 = sum__19[8] ? result_exp__59 : result_exp__60;
  assign x_bexp__820 = 8'h00;
  assign result_fraction__231 = is_result_nan__77 ? nan_fraction__131 : result_fraction__229;
  assign result_fraction__230 = is_result_nan__76 ? nan_fraction__130 : result_fraction__228;
  assign y_sq_bexp__6 = sum__38[8] ? result_exp__119 : result_exp__120;
  assign x_bexp__821 = 8'h00;
  assign result_fraction__348 = is_result_nan__116 ? nan_fraction__160 : result_fraction__346;
  assign result_fraction__347 = is_result_nan__115 ? nan_fraction__159 : result_fraction__345;
  assign y_sq_bexp__10 = sum__57[8] ? result_exp__179 : result_exp__180;
  assign x_bexp__822 = 8'h00;
  assign result_fraction__465 = is_result_nan__155 ? nan_fraction__189 : result_fraction__463;
  assign result_fraction__464 = is_result_nan__154 ? nan_fraction__188 : result_fraction__462;
  assign y_sq_bexp__14 = sum__76[8] ? result_exp__239 : result_exp__240;
  assign x_bexp__823 = 8'h00;
  assign y_sq_fraction = sum__19[8] ? result_fraction__113 : result_fraction__114;
  assign incremented_sum__94 = sum__19[7:0] + 8'h01;
  assign y_sq_fraction__3 = sum__38[8] ? result_fraction__230 : result_fraction__231;
  assign incremented_sum__112 = sum__38[7:0] + 8'h01;
  assign y_sq_fraction__6 = sum__57[8] ? result_fraction__347 : result_fraction__348;
  assign incremented_sum__130 = sum__57[7:0] + 8'h01;
  assign y_sq_fraction__9 = sum__76[8] ? result_fraction__464 : result_fraction__465;
  assign incremented_sum__148 = sum__76[7:0] + 8'h01;
  assign wide_y__37 = {2'h1, y_sq_fraction, 3'h0};
  assign x_sq_bexpbs_difference__1 = sum__19[8] ? incremented_sum__94 : ~sum__19[7:0];
  assign wide_y__75 = {2'h1, y_sq_fraction__3, 3'h0};
  assign x_sq_bexpbs_difference__2 = sum__38[8] ? incremented_sum__112 : ~sum__38[7:0];
  assign wide_y__113 = {2'h1, y_sq_fraction__6, 3'h0};
  assign x_sq_bexpbs_difference__3 = sum__57[8] ? incremented_sum__130 : ~sum__57[7:0];
  assign wide_y__151 = {2'h1, y_sq_fraction__9, 3'h0};
  assign x_sq_bexpbs_difference__4 = sum__76[8] ? incremented_sum__148 : ~sum__76[7:0];
  assign wide_y__38 = wide_y__37 & {28{y_sq_bexp__1 != x_bexp__820}};
  assign sub_172687 = 8'h1c - x_sq_bexpbs_difference__1;
  assign wide_y__76 = wide_y__75 & {28{y_sq_bexp__6 != x_bexp__821}};
  assign sub_172689 = 8'h1c - x_sq_bexpbs_difference__2;
  assign wide_y__114 = wide_y__113 & {28{y_sq_bexp__10 != x_bexp__822}};
  assign sub_172691 = 8'h1c - x_sq_bexpbs_difference__3;
  assign wide_y__152 = wide_y__151 & {28{y_sq_bexp__14 != x_bexp__823}};
  assign sub_172693 = 8'h1c - x_sq_bexpbs_difference__4;
  assign dropped__19 = sub_172687 >= 8'h1c ? 28'h000_0000 : wide_y__38 << sub_172687;
  assign dropped__38 = sub_172689 >= 8'h1c ? 28'h000_0000 : wide_y__76 << sub_172689;
  assign dropped__57 = sub_172691 >= 8'h1c ? 28'h000_0000 : wide_y__114 << sub_172691;
  assign dropped__76 = sub_172693 >= 8'h1c ? 28'h000_0000 : wide_y__152 << sub_172693;
  assign x_sq_bexp__2 = sum__19[8] ? result_exp__60 : result_exp__59;
  assign x_bexp__824 = 8'h00;
  assign x_sq_bexp__5 = sum__38[8] ? result_exp__120 : result_exp__119;
  assign x_bexp__825 = 8'h00;
  assign x_sq_bexp__10 = sum__57[8] ? result_exp__180 : result_exp__179;
  assign x_bexp__826 = 8'h00;
  assign x_sq_bexp__14 = sum__76[8] ? result_exp__240 : result_exp__239;
  assign x_bexp__827 = 8'h00;
  assign x_sq_fraction = sum__19[8] ? result_fraction__114 : result_fraction__113;
  assign sticky__59 = {27'h000_0000, dropped__19[27:3] != 25'h000_0000};
  assign x_sq_fraction__1 = sum__38[8] ? result_fraction__231 : result_fraction__230;
  assign sticky__118 = {27'h000_0000, dropped__38[27:3] != 25'h000_0000};
  assign x_sq_fraction__6 = sum__57[8] ? result_fraction__348 : result_fraction__347;
  assign sticky__177 = {27'h000_0000, dropped__57[27:3] != 25'h000_0000};
  assign x_sq_fraction__9 = sum__76[8] ? result_fraction__465 : result_fraction__464;
  assign sticky__236 = {27'h000_0000, dropped__76[27:3] != 25'h000_0000};
  assign x_sqddend_y = (x_sq_bexpbs_difference__1 >= 8'h1c ? 28'h000_0000 : wide_y__38 >> x_sq_bexpbs_difference__1) | sticky__59;
  assign x_sqddend_y__1 = (x_sq_bexpbs_difference__2 >= 8'h1c ? 28'h000_0000 : wide_y__76 >> x_sq_bexpbs_difference__2) | sticky__118;
  assign x_sqddend_y__2 = (x_sq_bexpbs_difference__3 >= 8'h1c ? 28'h000_0000 : wide_y__114 >> x_sq_bexpbs_difference__3) | sticky__177;
  assign x_sqddend_y__3 = (x_sq_bexpbs_difference__4 >= 8'h1c ? 28'h000_0000 : wide_y__152 >> x_sq_bexpbs_difference__4) | sticky__236;
  assign wide_x__153 = {2'h1, x_sq_fraction} & {25{x_sq_bexp__2 != x_bexp__824}};
  assign wide_x__154 = {2'h1, x_sq_fraction__1} & {25{x_sq_bexp__5 != x_bexp__825}};
  assign wide_x__155 = {2'h1, x_sq_fraction__6} & {25{x_sq_bexp__10 != x_bexp__826}};
  assign wide_x__156 = {2'h1, x_sq_fraction__9} & {25{x_sq_bexp__14 != x_bexp__827}};
  assign bit_slice_172762 = x_sqddend_y[2:0];
  assign carry_fraction__155 = wide_x__153 + x_sqddend_y[27:3];
  assign bit_slice_172764 = x_sqddend_y__1[2:0];
  assign carry_fraction__158 = wide_x__154 + x_sqddend_y__1[27:3];
  assign bit_slice_172766 = x_sqddend_y__2[2:0];
  assign carry_fraction__161 = wide_x__155 + x_sqddend_y__2[27:3];
  assign bit_slice_172768 = x_sqddend_y__3[2:0];
  assign carry_fraction__164 = wide_x__156 + x_sqddend_y__3[27:3];
  assign concat_172778 = {{bit_slice_172762[0], bit_slice_172762[1], bit_slice_172762[2]}, {carry_fraction__155[0], carry_fraction__155[1], carry_fraction__155[2], carry_fraction__155[3], carry_fraction__155[4], carry_fraction__155[5], carry_fraction__155[6], carry_fraction__155[7], carry_fraction__155[8], carry_fraction__155[9], carry_fraction__155[10], carry_fraction__155[11], carry_fraction__155[12], carry_fraction__155[13], carry_fraction__155[14], carry_fraction__155[15], carry_fraction__155[16], carry_fraction__155[17], carry_fraction__155[18], carry_fraction__155[19], carry_fraction__155[20], carry_fraction__155[21], carry_fraction__155[22], carry_fraction__155[23], carry_fraction__155[24]}};
  assign concat_172779 = {{bit_slice_172764[0], bit_slice_172764[1], bit_slice_172764[2]}, {carry_fraction__158[0], carry_fraction__158[1], carry_fraction__158[2], carry_fraction__158[3], carry_fraction__158[4], carry_fraction__158[5], carry_fraction__158[6], carry_fraction__158[7], carry_fraction__158[8], carry_fraction__158[9], carry_fraction__158[10], carry_fraction__158[11], carry_fraction__158[12], carry_fraction__158[13], carry_fraction__158[14], carry_fraction__158[15], carry_fraction__158[16], carry_fraction__158[17], carry_fraction__158[18], carry_fraction__158[19], carry_fraction__158[20], carry_fraction__158[21], carry_fraction__158[22], carry_fraction__158[23], carry_fraction__158[24]}};
  assign concat_172780 = {{bit_slice_172766[0], bit_slice_172766[1], bit_slice_172766[2]}, {carry_fraction__161[0], carry_fraction__161[1], carry_fraction__161[2], carry_fraction__161[3], carry_fraction__161[4], carry_fraction__161[5], carry_fraction__161[6], carry_fraction__161[7], carry_fraction__161[8], carry_fraction__161[9], carry_fraction__161[10], carry_fraction__161[11], carry_fraction__161[12], carry_fraction__161[13], carry_fraction__161[14], carry_fraction__161[15], carry_fraction__161[16], carry_fraction__161[17], carry_fraction__161[18], carry_fraction__161[19], carry_fraction__161[20], carry_fraction__161[21], carry_fraction__161[22], carry_fraction__161[23], carry_fraction__161[24]}};
  assign concat_172781 = {{bit_slice_172768[0], bit_slice_172768[1], bit_slice_172768[2]}, {carry_fraction__164[0], carry_fraction__164[1], carry_fraction__164[2], carry_fraction__164[3], carry_fraction__164[4], carry_fraction__164[5], carry_fraction__164[6], carry_fraction__164[7], carry_fraction__164[8], carry_fraction__164[9], carry_fraction__164[10], carry_fraction__164[11], carry_fraction__164[12], carry_fraction__164[13], carry_fraction__164[14], carry_fraction__164[15], carry_fraction__164[16], carry_fraction__164[17], carry_fraction__164[18], carry_fraction__164[19], carry_fraction__164[20], carry_fraction__164[21], carry_fraction__164[22], carry_fraction__164[23], carry_fraction__164[24]}};
  assign one_hot_172782 = {concat_172778[27:0] == 28'h000_0000, concat_172778[27] && concat_172778[26:0] == 27'h000_0000, concat_172778[26] && concat_172778[25:0] == 26'h000_0000, concat_172778[25] && concat_172778[24:0] == 25'h000_0000, concat_172778[24] && concat_172778[23:0] == 24'h00_0000, concat_172778[23] && concat_172778[22:0] == 23'h00_0000, concat_172778[22] && concat_172778[21:0] == 22'h00_0000, concat_172778[21] && concat_172778[20:0] == 21'h00_0000, concat_172778[20] && concat_172778[19:0] == 20'h0_0000, concat_172778[19] && concat_172778[18:0] == 19'h0_0000, concat_172778[18] && concat_172778[17:0] == 18'h0_0000, concat_172778[17] && concat_172778[16:0] == 17'h0_0000, concat_172778[16] && concat_172778[15:0] == 16'h0000, concat_172778[15] && concat_172778[14:0] == 15'h0000, concat_172778[14] && concat_172778[13:0] == 14'h0000, concat_172778[13] && concat_172778[12:0] == 13'h0000, concat_172778[12] && concat_172778[11:0] == 12'h000, concat_172778[11] && concat_172778[10:0] == 11'h000, concat_172778[10] && concat_172778[9:0] == 10'h000, concat_172778[9] && concat_172778[8:0] == 9'h000, concat_172778[8] && concat_172778[7:0] == 8'h00, concat_172778[7] && concat_172778[6:0] == 7'h00, concat_172778[6] && concat_172778[5:0] == 6'h00, concat_172778[5] && concat_172778[4:0] == 5'h00, concat_172778[4] && concat_172778[3:0] == 4'h0, concat_172778[3] && concat_172778[2:0] == 3'h0, concat_172778[2] && concat_172778[1:0] == 2'h0, concat_172778[1] && !concat_172778[0], concat_172778[0]};
  assign one_hot_172783 = {concat_172779[27:0] == 28'h000_0000, concat_172779[27] && concat_172779[26:0] == 27'h000_0000, concat_172779[26] && concat_172779[25:0] == 26'h000_0000, concat_172779[25] && concat_172779[24:0] == 25'h000_0000, concat_172779[24] && concat_172779[23:0] == 24'h00_0000, concat_172779[23] && concat_172779[22:0] == 23'h00_0000, concat_172779[22] && concat_172779[21:0] == 22'h00_0000, concat_172779[21] && concat_172779[20:0] == 21'h00_0000, concat_172779[20] && concat_172779[19:0] == 20'h0_0000, concat_172779[19] && concat_172779[18:0] == 19'h0_0000, concat_172779[18] && concat_172779[17:0] == 18'h0_0000, concat_172779[17] && concat_172779[16:0] == 17'h0_0000, concat_172779[16] && concat_172779[15:0] == 16'h0000, concat_172779[15] && concat_172779[14:0] == 15'h0000, concat_172779[14] && concat_172779[13:0] == 14'h0000, concat_172779[13] && concat_172779[12:0] == 13'h0000, concat_172779[12] && concat_172779[11:0] == 12'h000, concat_172779[11] && concat_172779[10:0] == 11'h000, concat_172779[10] && concat_172779[9:0] == 10'h000, concat_172779[9] && concat_172779[8:0] == 9'h000, concat_172779[8] && concat_172779[7:0] == 8'h00, concat_172779[7] && concat_172779[6:0] == 7'h00, concat_172779[6] && concat_172779[5:0] == 6'h00, concat_172779[5] && concat_172779[4:0] == 5'h00, concat_172779[4] && concat_172779[3:0] == 4'h0, concat_172779[3] && concat_172779[2:0] == 3'h0, concat_172779[2] && concat_172779[1:0] == 2'h0, concat_172779[1] && !concat_172779[0], concat_172779[0]};
  assign one_hot_172784 = {concat_172780[27:0] == 28'h000_0000, concat_172780[27] && concat_172780[26:0] == 27'h000_0000, concat_172780[26] && concat_172780[25:0] == 26'h000_0000, concat_172780[25] && concat_172780[24:0] == 25'h000_0000, concat_172780[24] && concat_172780[23:0] == 24'h00_0000, concat_172780[23] && concat_172780[22:0] == 23'h00_0000, concat_172780[22] && concat_172780[21:0] == 22'h00_0000, concat_172780[21] && concat_172780[20:0] == 21'h00_0000, concat_172780[20] && concat_172780[19:0] == 20'h0_0000, concat_172780[19] && concat_172780[18:0] == 19'h0_0000, concat_172780[18] && concat_172780[17:0] == 18'h0_0000, concat_172780[17] && concat_172780[16:0] == 17'h0_0000, concat_172780[16] && concat_172780[15:0] == 16'h0000, concat_172780[15] && concat_172780[14:0] == 15'h0000, concat_172780[14] && concat_172780[13:0] == 14'h0000, concat_172780[13] && concat_172780[12:0] == 13'h0000, concat_172780[12] && concat_172780[11:0] == 12'h000, concat_172780[11] && concat_172780[10:0] == 11'h000, concat_172780[10] && concat_172780[9:0] == 10'h000, concat_172780[9] && concat_172780[8:0] == 9'h000, concat_172780[8] && concat_172780[7:0] == 8'h00, concat_172780[7] && concat_172780[6:0] == 7'h00, concat_172780[6] && concat_172780[5:0] == 6'h00, concat_172780[5] && concat_172780[4:0] == 5'h00, concat_172780[4] && concat_172780[3:0] == 4'h0, concat_172780[3] && concat_172780[2:0] == 3'h0, concat_172780[2] && concat_172780[1:0] == 2'h0, concat_172780[1] && !concat_172780[0], concat_172780[0]};
  assign one_hot_172785 = {concat_172781[27:0] == 28'h000_0000, concat_172781[27] && concat_172781[26:0] == 27'h000_0000, concat_172781[26] && concat_172781[25:0] == 26'h000_0000, concat_172781[25] && concat_172781[24:0] == 25'h000_0000, concat_172781[24] && concat_172781[23:0] == 24'h00_0000, concat_172781[23] && concat_172781[22:0] == 23'h00_0000, concat_172781[22] && concat_172781[21:0] == 22'h00_0000, concat_172781[21] && concat_172781[20:0] == 21'h00_0000, concat_172781[20] && concat_172781[19:0] == 20'h0_0000, concat_172781[19] && concat_172781[18:0] == 19'h0_0000, concat_172781[18] && concat_172781[17:0] == 18'h0_0000, concat_172781[17] && concat_172781[16:0] == 17'h0_0000, concat_172781[16] && concat_172781[15:0] == 16'h0000, concat_172781[15] && concat_172781[14:0] == 15'h0000, concat_172781[14] && concat_172781[13:0] == 14'h0000, concat_172781[13] && concat_172781[12:0] == 13'h0000, concat_172781[12] && concat_172781[11:0] == 12'h000, concat_172781[11] && concat_172781[10:0] == 11'h000, concat_172781[10] && concat_172781[9:0] == 10'h000, concat_172781[9] && concat_172781[8:0] == 9'h000, concat_172781[8] && concat_172781[7:0] == 8'h00, concat_172781[7] && concat_172781[6:0] == 7'h00, concat_172781[6] && concat_172781[5:0] == 6'h00, concat_172781[5] && concat_172781[4:0] == 5'h00, concat_172781[4] && concat_172781[3:0] == 4'h0, concat_172781[3] && concat_172781[2:0] == 3'h0, concat_172781[2] && concat_172781[1:0] == 2'h0, concat_172781[1] && !concat_172781[0], concat_172781[0]};
  assign encode_172786 = {one_hot_172782[16] | one_hot_172782[17] | one_hot_172782[18] | one_hot_172782[19] | one_hot_172782[20] | one_hot_172782[21] | one_hot_172782[22] | one_hot_172782[23] | one_hot_172782[24] | one_hot_172782[25] | one_hot_172782[26] | one_hot_172782[27] | one_hot_172782[28], one_hot_172782[8] | one_hot_172782[9] | one_hot_172782[10] | one_hot_172782[11] | one_hot_172782[12] | one_hot_172782[13] | one_hot_172782[14] | one_hot_172782[15] | one_hot_172782[24] | one_hot_172782[25] | one_hot_172782[26] | one_hot_172782[27] | one_hot_172782[28], one_hot_172782[4] | one_hot_172782[5] | one_hot_172782[6] | one_hot_172782[7] | one_hot_172782[12] | one_hot_172782[13] | one_hot_172782[14] | one_hot_172782[15] | one_hot_172782[20] | one_hot_172782[21] | one_hot_172782[22] | one_hot_172782[23] | one_hot_172782[28], one_hot_172782[2] | one_hot_172782[3] | one_hot_172782[6] | one_hot_172782[7] | one_hot_172782[10] | one_hot_172782[11] | one_hot_172782[14] | one_hot_172782[15] | one_hot_172782[18] | one_hot_172782[19] | one_hot_172782[22] | one_hot_172782[23] | one_hot_172782[26] | one_hot_172782[27], one_hot_172782[1] | one_hot_172782[3] | one_hot_172782[5] | one_hot_172782[7] | one_hot_172782[9] | one_hot_172782[11] | one_hot_172782[13] | one_hot_172782[15] | one_hot_172782[17] | one_hot_172782[19] | one_hot_172782[21] | one_hot_172782[23] | one_hot_172782[25] | one_hot_172782[27]};
  assign encode_172787 = {one_hot_172783[16] | one_hot_172783[17] | one_hot_172783[18] | one_hot_172783[19] | one_hot_172783[20] | one_hot_172783[21] | one_hot_172783[22] | one_hot_172783[23] | one_hot_172783[24] | one_hot_172783[25] | one_hot_172783[26] | one_hot_172783[27] | one_hot_172783[28], one_hot_172783[8] | one_hot_172783[9] | one_hot_172783[10] | one_hot_172783[11] | one_hot_172783[12] | one_hot_172783[13] | one_hot_172783[14] | one_hot_172783[15] | one_hot_172783[24] | one_hot_172783[25] | one_hot_172783[26] | one_hot_172783[27] | one_hot_172783[28], one_hot_172783[4] | one_hot_172783[5] | one_hot_172783[6] | one_hot_172783[7] | one_hot_172783[12] | one_hot_172783[13] | one_hot_172783[14] | one_hot_172783[15] | one_hot_172783[20] | one_hot_172783[21] | one_hot_172783[22] | one_hot_172783[23] | one_hot_172783[28], one_hot_172783[2] | one_hot_172783[3] | one_hot_172783[6] | one_hot_172783[7] | one_hot_172783[10] | one_hot_172783[11] | one_hot_172783[14] | one_hot_172783[15] | one_hot_172783[18] | one_hot_172783[19] | one_hot_172783[22] | one_hot_172783[23] | one_hot_172783[26] | one_hot_172783[27], one_hot_172783[1] | one_hot_172783[3] | one_hot_172783[5] | one_hot_172783[7] | one_hot_172783[9] | one_hot_172783[11] | one_hot_172783[13] | one_hot_172783[15] | one_hot_172783[17] | one_hot_172783[19] | one_hot_172783[21] | one_hot_172783[23] | one_hot_172783[25] | one_hot_172783[27]};
  assign encode_172788 = {one_hot_172784[16] | one_hot_172784[17] | one_hot_172784[18] | one_hot_172784[19] | one_hot_172784[20] | one_hot_172784[21] | one_hot_172784[22] | one_hot_172784[23] | one_hot_172784[24] | one_hot_172784[25] | one_hot_172784[26] | one_hot_172784[27] | one_hot_172784[28], one_hot_172784[8] | one_hot_172784[9] | one_hot_172784[10] | one_hot_172784[11] | one_hot_172784[12] | one_hot_172784[13] | one_hot_172784[14] | one_hot_172784[15] | one_hot_172784[24] | one_hot_172784[25] | one_hot_172784[26] | one_hot_172784[27] | one_hot_172784[28], one_hot_172784[4] | one_hot_172784[5] | one_hot_172784[6] | one_hot_172784[7] | one_hot_172784[12] | one_hot_172784[13] | one_hot_172784[14] | one_hot_172784[15] | one_hot_172784[20] | one_hot_172784[21] | one_hot_172784[22] | one_hot_172784[23] | one_hot_172784[28], one_hot_172784[2] | one_hot_172784[3] | one_hot_172784[6] | one_hot_172784[7] | one_hot_172784[10] | one_hot_172784[11] | one_hot_172784[14] | one_hot_172784[15] | one_hot_172784[18] | one_hot_172784[19] | one_hot_172784[22] | one_hot_172784[23] | one_hot_172784[26] | one_hot_172784[27], one_hot_172784[1] | one_hot_172784[3] | one_hot_172784[5] | one_hot_172784[7] | one_hot_172784[9] | one_hot_172784[11] | one_hot_172784[13] | one_hot_172784[15] | one_hot_172784[17] | one_hot_172784[19] | one_hot_172784[21] | one_hot_172784[23] | one_hot_172784[25] | one_hot_172784[27]};
  assign encode_172789 = {one_hot_172785[16] | one_hot_172785[17] | one_hot_172785[18] | one_hot_172785[19] | one_hot_172785[20] | one_hot_172785[21] | one_hot_172785[22] | one_hot_172785[23] | one_hot_172785[24] | one_hot_172785[25] | one_hot_172785[26] | one_hot_172785[27] | one_hot_172785[28], one_hot_172785[8] | one_hot_172785[9] | one_hot_172785[10] | one_hot_172785[11] | one_hot_172785[12] | one_hot_172785[13] | one_hot_172785[14] | one_hot_172785[15] | one_hot_172785[24] | one_hot_172785[25] | one_hot_172785[26] | one_hot_172785[27] | one_hot_172785[28], one_hot_172785[4] | one_hot_172785[5] | one_hot_172785[6] | one_hot_172785[7] | one_hot_172785[12] | one_hot_172785[13] | one_hot_172785[14] | one_hot_172785[15] | one_hot_172785[20] | one_hot_172785[21] | one_hot_172785[22] | one_hot_172785[23] | one_hot_172785[28], one_hot_172785[2] | one_hot_172785[3] | one_hot_172785[6] | one_hot_172785[7] | one_hot_172785[10] | one_hot_172785[11] | one_hot_172785[14] | one_hot_172785[15] | one_hot_172785[18] | one_hot_172785[19] | one_hot_172785[22] | one_hot_172785[23] | one_hot_172785[26] | one_hot_172785[27], one_hot_172785[1] | one_hot_172785[3] | one_hot_172785[5] | one_hot_172785[7] | one_hot_172785[9] | one_hot_172785[11] | one_hot_172785[13] | one_hot_172785[15] | one_hot_172785[17] | one_hot_172785[19] | one_hot_172785[21] | one_hot_172785[23] | one_hot_172785[25] | one_hot_172785[27]};
  assign cancel__19 = |encode_172786[4:1];
  assign carry_bit__19 = carry_fraction__155[24];
  assign result_fraction__536 = 23'h00_0000;
  assign cancel__38 = |encode_172787[4:1];
  assign carry_bit__38 = carry_fraction__158[24];
  assign result_fraction__603 = 23'h00_0000;
  assign cancel__57 = |encode_172788[4:1];
  assign carry_bit__57 = carry_fraction__161[24];
  assign result_fraction__670 = 23'h00_0000;
  assign cancel__76 = |encode_172789[4:1];
  assign carry_bit__76 = carry_fraction__164[24];
  assign result_fraction__749 = 23'h00_0000;
  assign leading_zeroes__19 = {result_fraction__536, encode_172786};
  assign leading_zeroes__38 = {result_fraction__603, encode_172787};
  assign leading_zeroes__57 = {result_fraction__670, encode_172788};
  assign leading_zeroes__76 = {result_fraction__749, encode_172789};
  assign carry_fraction__154 = x_sqddend_y[2];
  assign carry_fraction__153 = x_sqddend_y[1] | x_sqddend_y[0];
  assign concat_172839 = {carry_fraction__155[23:0], bit_slice_172762};
  assign add_172840 = leading_zeroes__19 + 28'hfff_ffff;
  assign carry_fraction__157 = x_sqddend_y__1[2];
  assign carry_fraction__156 = x_sqddend_y__1[1] | x_sqddend_y__1[0];
  assign concat_172846 = {carry_fraction__158[23:0], bit_slice_172764};
  assign add_172847 = leading_zeroes__38 + 28'hfff_ffff;
  assign carry_fraction__160 = x_sqddend_y__2[2];
  assign carry_fraction__159 = x_sqddend_y__2[1] | x_sqddend_y__2[0];
  assign concat_172853 = {carry_fraction__161[23:0], bit_slice_172766};
  assign add_172854 = leading_zeroes__57 + 28'hfff_ffff;
  assign carry_fraction__163 = x_sqddend_y__3[2];
  assign carry_fraction__162 = x_sqddend_y__3[1] | x_sqddend_y__3[0];
  assign concat_172860 = {carry_fraction__164[23:0], bit_slice_172768};
  assign add_172861 = leading_zeroes__76 + 28'hfff_ffff;
  assign concat_172862 = {~(carry_bit__19 | cancel__19), ~(carry_bit__19 | ~cancel__19), ~(~carry_bit__19 | cancel__19)};
  assign carry_fraction__38 = {carry_fraction__155, carry_fraction__154, carry_fraction__153};
  assign cancel_fraction__19 = add_172840 >= 28'h000_001b ? 27'h000_0000 : concat_172839 << add_172840;
  assign concat_172865 = {~(carry_bit__38 | cancel__38), ~(carry_bit__38 | ~cancel__38), ~(~carry_bit__38 | cancel__38)};
  assign carry_fraction__76 = {carry_fraction__158, carry_fraction__157, carry_fraction__156};
  assign cancel_fraction__38 = add_172847 >= 28'h000_001b ? 27'h000_0000 : concat_172846 << add_172847;
  assign concat_172868 = {~(carry_bit__57 | cancel__57), ~(carry_bit__57 | ~cancel__57), ~(~carry_bit__57 | cancel__57)};
  assign carry_fraction__114 = {carry_fraction__161, carry_fraction__160, carry_fraction__159};
  assign cancel_fraction__57 = add_172854 >= 28'h000_001b ? 27'h000_0000 : concat_172853 << add_172854;
  assign concat_172871 = {~(carry_bit__76 | cancel__76), ~(carry_bit__76 | ~cancel__76), ~(~carry_bit__76 | cancel__76)};
  assign carry_fraction__152 = {carry_fraction__164, carry_fraction__163, carry_fraction__162};
  assign cancel_fraction__76 = add_172861 >= 28'h000_001b ? 27'h000_0000 : concat_172860 << add_172861;
  assign shifted_fraction__19 = carry_fraction__38 & {27{concat_172862[0]}} | cancel_fraction__19 & {27{concat_172862[1]}} | concat_172839 & {27{concat_172862[2]}};
  assign shifted_fraction__38 = carry_fraction__76 & {27{concat_172865[0]}} | cancel_fraction__38 & {27{concat_172865[1]}} | concat_172846 & {27{concat_172865[2]}};
  assign shifted_fraction__57 = carry_fraction__114 & {27{concat_172868[0]}} | cancel_fraction__57 & {27{concat_172868[1]}} | concat_172853 & {27{concat_172868[2]}};
  assign shifted_fraction__76 = carry_fraction__152 & {27{concat_172871[0]}} | cancel_fraction__76 & {27{concat_172871[1]}} | concat_172860 & {27{concat_172871[2]}};
  assign result_sign__1100 = 1'h0;
  assign result_sign__1101 = 1'h0;
  assign result_sign__1102 = 1'h0;
  assign result_sign__1103 = 1'h0;
  assign normal_chunk__19 = shifted_fraction__19[2:0];
  assign fraction_shift__261 = 3'h4;
  assign half_way_chunk__19 = shifted_fraction__19[3:2];
  assign normal_chunk__38 = shifted_fraction__38[2:0];
  assign fraction_shift__296 = 3'h4;
  assign half_way_chunk__38 = shifted_fraction__38[3:2];
  assign normal_chunk__57 = shifted_fraction__57[2:0];
  assign fraction_shift__331 = 3'h4;
  assign half_way_chunk__57 = shifted_fraction__57[3:2];
  assign normal_chunk__76 = shifted_fraction__76[2:0];
  assign fraction_shift__366 = 3'h4;
  assign half_way_chunk__76 = shifted_fraction__76[3:2];
  assign result_sign__478 = 1'h0;
  assign add_172913 = {result_sign__1100, shifted_fraction__19[26:3]} + 25'h000_0001;
  assign result_sign__575 = 1'h0;
  assign add_172917 = {result_sign__1101, shifted_fraction__38[26:3]} + 25'h000_0001;
  assign result_sign__677 = 1'h0;
  assign add_172921 = {result_sign__1102, shifted_fraction__57[26:3]} + 25'h000_0001;
  assign result_sign__789 = 1'h0;
  assign add_172925 = {result_sign__1103, shifted_fraction__76[26:3]} + 25'h000_0001;
  assign do_round_up__39 = normal_chunk__19 > fraction_shift__261 | half_way_chunk__19 == 2'h3;
  assign do_round_up__78 = normal_chunk__38 > fraction_shift__296 | half_way_chunk__38 == 2'h3;
  assign do_round_up__117 = normal_chunk__57 > fraction_shift__331 | half_way_chunk__57 == 2'h3;
  assign do_round_up__156 = normal_chunk__76 > fraction_shift__366 | half_way_chunk__76 == 2'h3;
  assign rounded_fraction__19 = do_round_up__39 ? {add_172913, normal_chunk__19} : {result_sign__478, shifted_fraction__19};
  assign rounded_fraction__38 = do_round_up__78 ? {add_172917, normal_chunk__38} : {result_sign__575, shifted_fraction__38};
  assign rounded_fraction__57 = do_round_up__117 ? {add_172921, normal_chunk__57} : {result_sign__677, shifted_fraction__57};
  assign rounded_fraction__76 = do_round_up__156 ? {add_172925, normal_chunk__76} : {result_sign__789, shifted_fraction__76};
  assign result_sign__479 = 1'h0;
  assign x_bexp__592 = 8'h00;
  assign rounding_carry__19 = rounded_fraction__19[27];
  assign result_sign__576 = 1'h0;
  assign x_bexp__610 = 8'h00;
  assign rounding_carry__38 = rounded_fraction__38[27];
  assign result_sign__678 = 1'h0;
  assign x_bexp__628 = 8'h00;
  assign rounding_carry__57 = rounded_fraction__57[27];
  assign result_sign__790 = 1'h0;
  assign x_bexp__646 = 8'h00;
  assign rounding_carry__76 = rounded_fraction__76[27];
  assign result_sign__480 = 1'h0;
  assign add_172963 = {result_sign__479, x_sq_bexp__2} + {x_bexp__592, rounding_carry__19};
  assign result_sign__577 = 1'h0;
  assign add_172967 = {result_sign__576, x_sq_bexp__5} + {x_bexp__610, rounding_carry__38};
  assign result_sign__679 = 1'h0;
  assign add_172971 = {result_sign__678, x_sq_bexp__10} + {x_bexp__628, rounding_carry__57};
  assign result_sign__791 = 1'h0;
  assign add_172975 = {result_sign__790, x_sq_bexp__14} + {x_bexp__646, rounding_carry__76};
  assign add_172998 = {result_sign__480, add_172963} + 10'h001;
  assign add_173001 = {result_sign__577, add_172967} + 10'h001;
  assign add_173004 = {result_sign__679, add_172971} + 10'h001;
  assign add_173007 = {result_sign__791, add_172975} + 10'h001;
  assign wide_exponent__55 = add_172998 - {5'h00, encode_172786};
  assign wide_exponent__112 = add_173001 - {5'h00, encode_172787};
  assign wide_exponent__169 = add_173004 - {5'h00, encode_172788};
  assign wide_exponent__226 = add_173007 - {5'h00, encode_172789};
  assign wide_exponent__56 = wide_exponent__55 & {10{carry_fraction__155 != 25'h000_0000 | bit_slice_172762 != 3'h0}};
  assign wide_exponent__113 = wide_exponent__112 & {10{carry_fraction__158 != 25'h000_0000 | bit_slice_172764 != 3'h0}};
  assign wide_exponent__170 = wide_exponent__169 & {10{carry_fraction__161 != 25'h000_0000 | bit_slice_172766 != 3'h0}};
  assign wide_exponent__227 = wide_exponent__226 & {10{carry_fraction__164 != 25'h000_0000 | bit_slice_172768 != 3'h0}};
  assign high_exp__138 = 8'hff;
  assign result_fraction__537 = 23'h00_0000;
  assign high_exp__139 = 8'hff;
  assign result_fraction__538 = 23'h00_0000;
  assign wide_exponent__57 = wide_exponent__56[8:0] & {9{~wide_exponent__56[9]}};
  assign high_exp__204 = 8'hff;
  assign result_fraction__604 = 23'h00_0000;
  assign high_exp__205 = 8'hff;
  assign result_fraction__605 = 23'h00_0000;
  assign wide_exponent__114 = wide_exponent__113[8:0] & {9{~wide_exponent__113[9]}};
  assign high_exp__272 = 8'hff;
  assign result_fraction__671 = 23'h00_0000;
  assign high_exp__273 = 8'hff;
  assign result_fraction__672 = 23'h00_0000;
  assign wide_exponent__171 = wide_exponent__170[8:0] & {9{~wide_exponent__170[9]}};
  assign high_exp__346 = 8'hff;
  assign result_fraction__750 = 23'h00_0000;
  assign high_exp__347 = 8'hff;
  assign result_fraction__751 = 23'h00_0000;
  assign wide_exponent__228 = wide_exponent__227[8:0] & {9{~wide_exponent__227[9]}};
  assign eq_173058 = x_sq_bexp__2 == high_exp__138;
  assign eq_173060 = y_sq_bexp__1 == high_exp__139;
  assign eq_173063 = x_sq_bexp__5 == high_exp__204;
  assign eq_173065 = y_sq_bexp__6 == high_exp__205;
  assign eq_173068 = x_sq_bexp__10 == high_exp__272;
  assign eq_173070 = y_sq_bexp__10 == high_exp__273;
  assign eq_173073 = x_sq_bexp__14 == high_exp__346;
  assign eq_173075 = y_sq_bexp__14 == high_exp__347;
  assign result_fraction__539 = 23'h00_0000;
  assign result_fraction__540 = 23'h00_0000;
  assign result_fraction__606 = 23'h00_0000;
  assign result_fraction__607 = 23'h00_0000;
  assign result_fraction__673 = 23'h00_0000;
  assign result_fraction__674 = 23'h00_0000;
  assign result_fraction__752 = 23'h00_0000;
  assign result_fraction__753 = 23'h00_0000;
  assign fraction_shift__384 = 3'h3;
  assign fraction_shift__262 = 3'h4;
  assign is_operand_inf__19 = eq_173058 & x_sq_fraction == result_fraction__537 | eq_173060 & y_sq_fraction == result_fraction__538;
  assign and_reduce_173112 = &wide_exponent__57[7:0];
  assign fraction_shift__402 = 3'h3;
  assign fraction_shift__297 = 3'h4;
  assign is_operand_inf__38 = eq_173063 & x_sq_fraction__1 == result_fraction__604 | eq_173065 & y_sq_fraction__3 == result_fraction__605;
  assign and_reduce_173120 = &wide_exponent__114[7:0];
  assign fraction_shift__420 = 3'h3;
  assign fraction_shift__332 = 3'h4;
  assign is_operand_inf__57 = eq_173068 & x_sq_fraction__6 == result_fraction__671 | eq_173070 & y_sq_fraction__6 == result_fraction__672;
  assign and_reduce_173128 = &wide_exponent__171[7:0];
  assign fraction_shift__438 = 3'h3;
  assign fraction_shift__367 = 3'h4;
  assign is_operand_inf__76 = eq_173073 & x_sq_fraction__9 == result_fraction__750 | eq_173075 & y_sq_fraction__9 == result_fraction__751;
  assign and_reduce_173136 = &wide_exponent__228[7:0];
  assign fraction_shift__57 = rounding_carry__19 ? fraction_shift__262 : fraction_shift__384;
  assign fraction_shift__114 = rounding_carry__38 ? fraction_shift__297 : fraction_shift__402;
  assign fraction_shift__171 = rounding_carry__57 ? fraction_shift__332 : fraction_shift__420;
  assign fraction_shift__228 = rounding_carry__76 ? fraction_shift__367 : fraction_shift__438;
  assign is_result_nan__39 = eq_173058 & x_sq_fraction != result_fraction__539 | eq_173060 & y_sq_fraction != result_fraction__540;
  assign shrl_173155 = rounded_fraction__19 >> fraction_shift__57;
  assign is_result_nan__78 = eq_173063 & x_sq_fraction__1 != result_fraction__606 | eq_173065 & y_sq_fraction__3 != result_fraction__607;
  assign shrl_173158 = rounded_fraction__38 >> fraction_shift__114;
  assign is_result_nan__117 = eq_173068 & x_sq_fraction__6 != result_fraction__673 | eq_173070 & y_sq_fraction__6 != result_fraction__674;
  assign shrl_173161 = rounded_fraction__57 >> fraction_shift__171;
  assign is_result_nan__156 = eq_173073 & x_sq_fraction__9 != result_fraction__752 | eq_173075 & y_sq_fraction__9 != result_fraction__753;
  assign shrl_173164 = rounded_fraction__76 >> fraction_shift__228;
  assign high_exp__140 = 8'hff;
  assign result_fraction__115 = shrl_173155[22:0];
  assign high_exp__206 = 8'hff;
  assign result_fraction__232 = shrl_173158[22:0];
  assign high_exp__274 = 8'hff;
  assign result_fraction__349 = shrl_173161[22:0];
  assign high_exp__348 = 8'hff;
  assign result_fraction__466 = shrl_173164[22:0];
  assign result_exponent__19 = is_result_nan__39 | is_operand_inf__19 | wide_exponent__57[8] | and_reduce_173112 ? high_exp__140 : wide_exponent__57[7:0];
  assign result_fraction__116 = result_fraction__115 & {23{~(is_operand_inf__19 | wide_exponent__57[8] | and_reduce_173112 | ~((|wide_exponent__57[8:1]) | wide_exponent__57[0]))}};
  assign nan_fraction__105 = 23'h40_0000;
  assign result_exponent__38 = is_result_nan__78 | is_operand_inf__38 | wide_exponent__114[8] | and_reduce_173120 ? high_exp__206 : wide_exponent__114[7:0];
  assign result_fraction__233 = result_fraction__232 & {23{~(is_operand_inf__38 | wide_exponent__114[8] | and_reduce_173120 | ~((|wide_exponent__114[8:1]) | wide_exponent__114[0]))}};
  assign nan_fraction__132 = 23'h40_0000;
  assign result_exponent__57 = is_result_nan__117 | is_operand_inf__57 | wide_exponent__171[8] | and_reduce_173128 ? high_exp__274 : wide_exponent__171[7:0];
  assign result_fraction__350 = result_fraction__349 & {23{~(is_operand_inf__57 | wide_exponent__171[8] | and_reduce_173128 | ~((|wide_exponent__171[8:1]) | wide_exponent__171[0]))}};
  assign nan_fraction__161 = 23'h40_0000;
  assign result_exponent__76 = is_result_nan__156 | is_operand_inf__76 | wide_exponent__228[8] | and_reduce_173136 ? high_exp__348 : wide_exponent__228[7:0];
  assign result_fraction__467 = result_fraction__466 & {23{~(is_operand_inf__76 | wide_exponent__228[8] | and_reduce_173136 | ~((|wide_exponent__228[8:1]) | wide_exponent__228[0]))}};
  assign nan_fraction__190 = 23'h40_0000;
  assign uexp = result_exponent__19 + 8'h81;
  assign result_fraction__117 = is_result_nan__39 ? nan_fraction__105 : result_fraction__116;
  assign result_sign__828 = 1'h0;
  assign uexp__1 = result_exponent__38 + 8'h81;
  assign result_fraction__234 = is_result_nan__78 ? nan_fraction__132 : result_fraction__233;
  assign result_sign__829 = 1'h0;
  assign uexp__2 = result_exponent__57 + 8'h81;
  assign result_fraction__351 = is_result_nan__117 ? nan_fraction__161 : result_fraction__350;
  assign result_sign__830 = 1'h0;
  assign uexp__3 = result_exponent__76 + 8'h81;
  assign result_fraction__468 = is_result_nan__156 ? nan_fraction__190 : result_fraction__467;
  assign result_sign__831 = 1'h0;
  assign sel_173230 = uexp[0] ? {1'h1, result_fraction__117, result_sign__828} : {2'h1, result_fraction__117};
  assign sel_173231 = uexp__1[0] ? {1'h1, result_fraction__234, result_sign__829} : {2'h1, result_fraction__234};
  assign sel_173232 = uexp__2[0] ? {1'h1, result_fraction__351, result_sign__830} : {2'h1, result_fraction__351};
  assign sel_173233 = uexp__3[0] ? {1'h1, result_fraction__468, result_sign__831} : {2'h1, result_fraction__468};
  assign add_173250 = {5'h00, sel_173230[24:23]} + 7'h7f;
  assign add_173251 = {5'h00, sel_173231[24:23]} + 7'h7f;
  assign add_173252 = {5'h00, sel_173232[24:23]} + 7'h7f;
  assign add_173253 = {5'h00, sel_173233[24:23]} + 7'h7f;
  assign add_173276 = {add_173250[5:0], sel_173230[22:21]} + 8'hfb;
  assign add_173280 = {add_173251[5:0], sel_173231[22:21]} + 8'hfb;
  assign add_173284 = {add_173252[5:0], sel_173232[22:21]} + 8'hfb;
  assign add_173288 = {add_173253[5:0], sel_173233[22:21]} + 8'hfb;
  assign ugt_173291 = {add_173250, sel_173230[22:0]} > 30'h009f_ffff;
  assign ugt_173296 = {add_173251, sel_173231[22:0]} > 30'h009f_ffff;
  assign ugt_173301 = {add_173252, sel_173232[22:0]} > 30'h009f_ffff;
  assign ugt_173306 = {add_173253, sel_173233[22:0]} > 30'h009f_ffff;
  assign shifting_bit_mask__1 = 32'h0040_0000;
  assign sel_173312 = ugt_173291 ? {add_173276, sel_173230[20:0]} : {add_173250[5:0], sel_173230[22:0]};
  assign shifting_bit_mask__100 = 32'h0040_0000;
  assign sel_173315 = ugt_173296 ? {add_173280, sel_173231[20:0]} : {add_173251[5:0], sel_173231[22:0]};
  assign shifting_bit_mask__101 = 32'h0040_0000;
  assign sel_173318 = ugt_173301 ? {add_173284, sel_173232[20:0]} : {add_173252[5:0], sel_173232[22:0]};
  assign shifting_bit_mask__102 = 32'h0040_0000;
  assign sel_173321 = ugt_173306 ? {add_173288, sel_173233[20:0]} : {add_173253[5:0], sel_173233[22:0]};
  assign temp__2 = {7'h01, ugt_173291, 24'h00_0000} | shifting_bit_mask__1;
  assign result_sign__832 = 1'h0;
  assign temp__27 = {7'h01, ugt_173296, 24'h00_0000} | shifting_bit_mask__100;
  assign result_sign__833 = 1'h0;
  assign temp__52 = {7'h01, ugt_173301, 24'h00_0000} | shifting_bit_mask__101;
  assign result_sign__834 = 1'h0;
  assign temp__77 = {7'h01, ugt_173306, 24'h00_0000} | shifting_bit_mask__102;
  assign result_sign__835 = 1'h0;
  assign concat_173339 = {ugt_173291, result_sign__832};
  assign concat_173344 = {ugt_173296, result_sign__833};
  assign concat_173349 = {ugt_173301, result_sign__834};
  assign concat_173354 = {ugt_173306, result_sign__835};
  assign ule_173358 = temp__2[31:3] <= sel_173312;
  assign sub_173360 = {sel_173312[27:0], 3'h0} - temp__2[30:0];
  assign ule_173361 = temp__27[31:3] <= sel_173315;
  assign sub_173363 = {sel_173315[27:0], 3'h0} - temp__27[30:0];
  assign ule_173364 = temp__52[31:3] <= sel_173318;
  assign sub_173366 = {sel_173318[27:0], 3'h0} - temp__52[30:0];
  assign ule_173367 = temp__77[31:3] <= sel_173321;
  assign sub_173369 = {sel_173321[27:0], 3'h0} - temp__77[30:0];
  assign sel_173371 = ule_173358 ? concat_173339 | 2'h1 : concat_173339;
  assign result_fraction__888 = 23'h00_0000;
  assign sel_173375 = ule_173361 ? concat_173344 | 2'h1 : concat_173344;
  assign result_fraction__889 = 23'h00_0000;
  assign sel_173379 = ule_173364 ? concat_173349 | 2'h1 : concat_173349;
  assign result_fraction__890 = 23'h00_0000;
  assign sel_173383 = ule_173367 ? concat_173354 | 2'h1 : concat_173354;
  assign result_fraction__891 = 23'h00_0000;
  assign shifting_bit_mask__2 = 32'h0020_0000;
  assign sel_173388 = ule_173358 ? sub_173360[30:3] : sel_173312[27:0];
  assign shifting_bit_mask__103 = 32'h0020_0000;
  assign sel_173391 = ule_173361 ? sub_173363[30:3] : sel_173315[27:0];
  assign shifting_bit_mask__104 = 32'h0020_0000;
  assign sel_173394 = ule_173364 ? sub_173366[30:3] : sel_173318[27:0];
  assign shifting_bit_mask__105 = 32'h0020_0000;
  assign sel_173397 = ule_173367 ? sub_173369[30:3] : sel_173321[27:0];
  assign temp__3 = {7'h01, sel_173371, result_fraction__888} | shifting_bit_mask__2;
  assign result_sign__836 = 1'h0;
  assign temp__28 = {7'h01, sel_173375, result_fraction__889} | shifting_bit_mask__103;
  assign result_sign__837 = 1'h0;
  assign temp__53 = {7'h01, sel_173379, result_fraction__890} | shifting_bit_mask__104;
  assign result_sign__838 = 1'h0;
  assign temp__78 = {7'h01, sel_173383, result_fraction__891} | shifting_bit_mask__105;
  assign result_sign__839 = 1'h0;
  assign concat_173415 = {sel_173371, result_sign__836};
  assign concat_173420 = {sel_173375, result_sign__837};
  assign concat_173425 = {sel_173379, result_sign__838};
  assign concat_173430 = {sel_173383, result_sign__839};
  assign ule_173434 = temp__3[31:4] <= sel_173388;
  assign sub_173436 = {sel_173388[26:0], 4'h0} - temp__3[30:0];
  assign ule_173437 = temp__28[31:4] <= sel_173391;
  assign sub_173439 = {sel_173391[26:0], 4'h0} - temp__28[30:0];
  assign ule_173440 = temp__53[31:4] <= sel_173394;
  assign sub_173442 = {sel_173394[26:0], 4'h0} - temp__53[30:0];
  assign ule_173443 = temp__78[31:4] <= sel_173397;
  assign sub_173445 = {sel_173397[26:0], 4'h0} - temp__78[30:0];
  assign sel_173447 = ule_173434 ? concat_173415 | 3'h1 : concat_173415;
  assign sel_173451 = ule_173437 ? concat_173420 | 3'h1 : concat_173420;
  assign sel_173455 = ule_173440 ? concat_173425 | 3'h1 : concat_173425;
  assign sel_173459 = ule_173443 ? concat_173430 | 3'h1 : concat_173430;
  assign shifting_bit_mask__3 = 32'h0010_0000;
  assign sel_173464 = ule_173434 ? sub_173436[30:4] : sel_173388[26:0];
  assign shifting_bit_mask__106 = 32'h0010_0000;
  assign sel_173467 = ule_173437 ? sub_173439[30:4] : sel_173391[26:0];
  assign shifting_bit_mask__107 = 32'h0010_0000;
  assign sel_173470 = ule_173440 ? sub_173442[30:4] : sel_173394[26:0];
  assign shifting_bit_mask__108 = 32'h0010_0000;
  assign sel_173473 = ule_173443 ? sub_173445[30:4] : sel_173397[26:0];
  assign temp__4 = {7'h01, sel_173447, 22'h00_0000} | shifting_bit_mask__3;
  assign result_sign__840 = 1'h0;
  assign temp__29 = {7'h01, sel_173451, 22'h00_0000} | shifting_bit_mask__106;
  assign result_sign__841 = 1'h0;
  assign temp__54 = {7'h01, sel_173455, 22'h00_0000} | shifting_bit_mask__107;
  assign result_sign__842 = 1'h0;
  assign temp__79 = {7'h01, sel_173459, 22'h00_0000} | shifting_bit_mask__108;
  assign result_sign__843 = 1'h0;
  assign concat_173491 = {sel_173447, result_sign__840};
  assign concat_173496 = {sel_173451, result_sign__841};
  assign concat_173501 = {sel_173455, result_sign__842};
  assign concat_173506 = {sel_173459, result_sign__843};
  assign ule_173510 = temp__4[31:5] <= sel_173464;
  assign sub_173512 = {sel_173464[25:0], 5'h00} - temp__4[30:0];
  assign ule_173513 = temp__29[31:5] <= sel_173467;
  assign sub_173515 = {sel_173467[25:0], 5'h00} - temp__29[30:0];
  assign ule_173516 = temp__54[31:5] <= sel_173470;
  assign sub_173518 = {sel_173470[25:0], 5'h00} - temp__54[30:0];
  assign ule_173519 = temp__79[31:5] <= sel_173473;
  assign sub_173521 = {sel_173473[25:0], 5'h00} - temp__79[30:0];
  assign sel_173523 = ule_173510 ? concat_173491 | 4'h1 : concat_173491;
  assign sel_173527 = ule_173513 ? concat_173496 | 4'h1 : concat_173496;
  assign sel_173531 = ule_173516 ? concat_173501 | 4'h1 : concat_173501;
  assign sel_173535 = ule_173519 ? concat_173506 | 4'h1 : concat_173506;
  assign shifting_bit_mask__4 = 32'h0008_0000;
  assign sel_173540 = ule_173510 ? sub_173512[30:5] : sel_173464[25:0];
  assign shifting_bit_mask__109 = 32'h0008_0000;
  assign sel_173543 = ule_173513 ? sub_173515[30:5] : sel_173467[25:0];
  assign shifting_bit_mask__110 = 32'h0008_0000;
  assign sel_173546 = ule_173516 ? sub_173518[30:5] : sel_173470[25:0];
  assign shifting_bit_mask__111 = 32'h0008_0000;
  assign sel_173549 = ule_173519 ? sub_173521[30:5] : sel_173473[25:0];
  assign temp__5 = {7'h01, sel_173523, 21'h00_0000} | shifting_bit_mask__4;
  assign result_sign__844 = 1'h0;
  assign temp__30 = {7'h01, sel_173527, 21'h00_0000} | shifting_bit_mask__109;
  assign result_sign__845 = 1'h0;
  assign temp__55 = {7'h01, sel_173531, 21'h00_0000} | shifting_bit_mask__110;
  assign result_sign__846 = 1'h0;
  assign temp__80 = {7'h01, sel_173535, 21'h00_0000} | shifting_bit_mask__111;
  assign result_sign__847 = 1'h0;
  assign concat_173567 = {sel_173523, result_sign__844};
  assign concat_173572 = {sel_173527, result_sign__845};
  assign concat_173577 = {sel_173531, result_sign__846};
  assign concat_173582 = {sel_173535, result_sign__847};
  assign ule_173586 = temp__5[31:6] <= sel_173540;
  assign sub_173588 = {sel_173540[24:0], 6'h00} - temp__5[30:0];
  assign ule_173589 = temp__30[31:6] <= sel_173543;
  assign sub_173591 = {sel_173543[24:0], 6'h00} - temp__30[30:0];
  assign ule_173592 = temp__55[31:6] <= sel_173546;
  assign sub_173594 = {sel_173546[24:0], 6'h00} - temp__55[30:0];
  assign ule_173595 = temp__80[31:6] <= sel_173549;
  assign sub_173597 = {sel_173549[24:0], 6'h00} - temp__80[30:0];
  assign sel_173599 = ule_173586 ? concat_173567 | 5'h01 : concat_173567;
  assign sel_173603 = ule_173589 ? concat_173572 | 5'h01 : concat_173572;
  assign sel_173607 = ule_173592 ? concat_173577 | 5'h01 : concat_173577;
  assign sel_173611 = ule_173595 ? concat_173582 | 5'h01 : concat_173582;
  assign shifting_bit_mask__5 = 32'h0004_0000;
  assign sel_173616 = ule_173586 ? sub_173588[30:6] : sel_173540[24:0];
  assign shifting_bit_mask__112 = 32'h0004_0000;
  assign sel_173619 = ule_173589 ? sub_173591[30:6] : sel_173543[24:0];
  assign shifting_bit_mask__113 = 32'h0004_0000;
  assign sel_173622 = ule_173592 ? sub_173594[30:6] : sel_173546[24:0];
  assign shifting_bit_mask__114 = 32'h0004_0000;
  assign sel_173625 = ule_173595 ? sub_173597[30:6] : sel_173549[24:0];
  assign temp__6 = {7'h01, sel_173599, 20'h0_0000} | shifting_bit_mask__5;
  assign result_sign__848 = 1'h0;
  assign temp__31 = {7'h01, sel_173603, 20'h0_0000} | shifting_bit_mask__112;
  assign result_sign__849 = 1'h0;
  assign temp__56 = {7'h01, sel_173607, 20'h0_0000} | shifting_bit_mask__113;
  assign result_sign__850 = 1'h0;
  assign temp__81 = {7'h01, sel_173611, 20'h0_0000} | shifting_bit_mask__114;
  assign result_sign__851 = 1'h0;
  assign concat_173643 = {sel_173599, result_sign__848};
  assign concat_173648 = {sel_173603, result_sign__849};
  assign concat_173653 = {sel_173607, result_sign__850};
  assign concat_173658 = {sel_173611, result_sign__851};
  assign ule_173662 = temp__6[31:7] <= sel_173616;
  assign sub_173664 = {sel_173616[23:0], 7'h00} - temp__6[30:0];
  assign ule_173665 = temp__31[31:7] <= sel_173619;
  assign sub_173667 = {sel_173619[23:0], 7'h00} - temp__31[30:0];
  assign ule_173668 = temp__56[31:7] <= sel_173622;
  assign sub_173670 = {sel_173622[23:0], 7'h00} - temp__56[30:0];
  assign ule_173671 = temp__81[31:7] <= sel_173625;
  assign sub_173673 = {sel_173625[23:0], 7'h00} - temp__81[30:0];
  assign sel_173675 = ule_173662 ? concat_173643 | 6'h01 : concat_173643;
  assign sel_173679 = ule_173665 ? concat_173648 | 6'h01 : concat_173648;
  assign sel_173683 = ule_173668 ? concat_173653 | 6'h01 : concat_173653;
  assign sel_173687 = ule_173671 ? concat_173658 | 6'h01 : concat_173658;
  assign shifting_bit_mask__6 = 32'h0002_0000;
  assign sel_173692 = ule_173662 ? sub_173664[30:7] : sel_173616[23:0];
  assign shifting_bit_mask__115 = 32'h0002_0000;
  assign sel_173695 = ule_173665 ? sub_173667[30:7] : sel_173619[23:0];
  assign shifting_bit_mask__116 = 32'h0002_0000;
  assign sel_173698 = ule_173668 ? sub_173670[30:7] : sel_173622[23:0];
  assign shifting_bit_mask__117 = 32'h0002_0000;
  assign sel_173701 = ule_173671 ? sub_173673[30:7] : sel_173625[23:0];
  assign temp__7 = {7'h01, sel_173675, 19'h0_0000} | shifting_bit_mask__6;
  assign result_sign__852 = 1'h0;
  assign x_bexp__656 = 8'h00;
  assign temp__32 = {7'h01, sel_173679, 19'h0_0000} | shifting_bit_mask__115;
  assign result_sign__853 = 1'h0;
  assign x_bexp__658 = 8'h00;
  assign temp__57 = {7'h01, sel_173683, 19'h0_0000} | shifting_bit_mask__116;
  assign result_sign__854 = 1'h0;
  assign x_bexp__660 = 8'h00;
  assign temp__82 = {7'h01, sel_173687, 19'h0_0000} | shifting_bit_mask__117;
  assign result_sign__855 = 1'h0;
  assign x_bexp__662 = 8'h00;
  assign concat_173719 = {sel_173675, result_sign__852};
  assign concat_173724 = {sel_173679, result_sign__853};
  assign concat_173729 = {sel_173683, result_sign__854};
  assign concat_173734 = {sel_173687, result_sign__855};
  assign ule_173738 = temp__7[31:8] <= sel_173692;
  assign sub_173740 = {sel_173692[22:0], x_bexp__656} - temp__7[30:0];
  assign ule_173741 = temp__32[31:8] <= sel_173695;
  assign sub_173743 = {sel_173695[22:0], x_bexp__658} - temp__32[30:0];
  assign ule_173744 = temp__57[31:8] <= sel_173698;
  assign sub_173746 = {sel_173698[22:0], x_bexp__660} - temp__57[30:0];
  assign ule_173747 = temp__82[31:8] <= sel_173701;
  assign sub_173749 = {sel_173701[22:0], x_bexp__662} - temp__82[30:0];
  assign sel_173751 = ule_173738 ? concat_173719 | 7'h01 : concat_173719;
  assign sel_173755 = ule_173741 ? concat_173724 | 7'h01 : concat_173724;
  assign sel_173759 = ule_173744 ? concat_173729 | 7'h01 : concat_173729;
  assign sel_173763 = ule_173747 ? concat_173734 | 7'h01 : concat_173734;
  assign shifting_bit_mask__7 = 32'h0001_0000;
  assign sel_173768 = ule_173738 ? sub_173740[30:8] : sel_173692[22:0];
  assign shifting_bit_mask__118 = 32'h0001_0000;
  assign sel_173771 = ule_173741 ? sub_173743[30:8] : sel_173695[22:0];
  assign shifting_bit_mask__119 = 32'h0001_0000;
  assign sel_173774 = ule_173744 ? sub_173746[30:8] : sel_173698[22:0];
  assign shifting_bit_mask__120 = 32'h0001_0000;
  assign sel_173777 = ule_173747 ? sub_173749[30:8] : sel_173701[22:0];
  assign temp__8 = {7'h01, sel_173751, 18'h0_0000} | shifting_bit_mask__7;
  assign result_sign__856 = 1'h0;
  assign temp__33 = {7'h01, sel_173755, 18'h0_0000} | shifting_bit_mask__118;
  assign result_sign__857 = 1'h0;
  assign temp__58 = {7'h01, sel_173759, 18'h0_0000} | shifting_bit_mask__119;
  assign result_sign__858 = 1'h0;
  assign temp__83 = {7'h01, sel_173763, 18'h0_0000} | shifting_bit_mask__120;
  assign result_sign__859 = 1'h0;
  assign concat_173795 = {sel_173751, result_sign__856};
  assign concat_173800 = {sel_173755, result_sign__857};
  assign concat_173805 = {sel_173759, result_sign__858};
  assign concat_173810 = {sel_173763, result_sign__859};
  assign ule_173814 = temp__8[31:9] <= sel_173768;
  assign sub_173816 = {sel_173768[21:0], 9'h000} - temp__8[30:0];
  assign ule_173817 = temp__33[31:9] <= sel_173771;
  assign sub_173819 = {sel_173771[21:0], 9'h000} - temp__33[30:0];
  assign ule_173820 = temp__58[31:9] <= sel_173774;
  assign sub_173822 = {sel_173774[21:0], 9'h000} - temp__58[30:0];
  assign ule_173823 = temp__83[31:9] <= sel_173777;
  assign sub_173825 = {sel_173777[21:0], 9'h000} - temp__83[30:0];
  assign sel_173827 = ule_173814 ? concat_173795 | 8'h01 : concat_173795;
  assign sel_173831 = ule_173817 ? concat_173800 | 8'h01 : concat_173800;
  assign sel_173835 = ule_173820 ? concat_173805 | 8'h01 : concat_173805;
  assign sel_173839 = ule_173823 ? concat_173810 | 8'h01 : concat_173810;
  assign shifting_bit_mask__8 = 32'h0000_8000;
  assign sel_173844 = ule_173814 ? sub_173816[30:9] : sel_173768[21:0];
  assign shifting_bit_mask__121 = 32'h0000_8000;
  assign sel_173847 = ule_173817 ? sub_173819[30:9] : sel_173771[21:0];
  assign shifting_bit_mask__122 = 32'h0000_8000;
  assign sel_173850 = ule_173820 ? sub_173822[30:9] : sel_173774[21:0];
  assign shifting_bit_mask__123 = 32'h0000_8000;
  assign sel_173853 = ule_173823 ? sub_173825[30:9] : sel_173777[21:0];
  assign temp__9 = {7'h01, sel_173827, 17'h0_0000} | shifting_bit_mask__8;
  assign result_sign__860 = 1'h0;
  assign temp__34 = {7'h01, sel_173831, 17'h0_0000} | shifting_bit_mask__121;
  assign result_sign__861 = 1'h0;
  assign temp__59 = {7'h01, sel_173835, 17'h0_0000} | shifting_bit_mask__122;
  assign result_sign__862 = 1'h0;
  assign temp__84 = {7'h01, sel_173839, 17'h0_0000} | shifting_bit_mask__123;
  assign result_sign__863 = 1'h0;
  assign concat_173871 = {sel_173827, result_sign__860};
  assign concat_173876 = {sel_173831, result_sign__861};
  assign concat_173881 = {sel_173835, result_sign__862};
  assign concat_173886 = {sel_173839, result_sign__863};
  assign ule_173890 = temp__9[31:10] <= sel_173844;
  assign sub_173892 = {sel_173844[20:0], 10'h000} - temp__9[30:0];
  assign ule_173893 = temp__34[31:10] <= sel_173847;
  assign sub_173895 = {sel_173847[20:0], 10'h000} - temp__34[30:0];
  assign ule_173896 = temp__59[31:10] <= sel_173850;
  assign sub_173898 = {sel_173850[20:0], 10'h000} - temp__59[30:0];
  assign ule_173899 = temp__84[31:10] <= sel_173853;
  assign sub_173901 = {sel_173853[20:0], 10'h000} - temp__84[30:0];
  assign sel_173903 = ule_173890 ? concat_173871 | 9'h001 : concat_173871;
  assign sel_173907 = ule_173893 ? concat_173876 | 9'h001 : concat_173876;
  assign sel_173911 = ule_173896 ? concat_173881 | 9'h001 : concat_173881;
  assign sel_173915 = ule_173899 ? concat_173886 | 9'h001 : concat_173886;
  assign shifting_bit_mask__9 = 32'h0000_4000;
  assign sel_173920 = ule_173890 ? sub_173892[30:10] : sel_173844[20:0];
  assign shifting_bit_mask__124 = 32'h0000_4000;
  assign sel_173923 = ule_173893 ? sub_173895[30:10] : sel_173847[20:0];
  assign shifting_bit_mask__125 = 32'h0000_4000;
  assign sel_173926 = ule_173896 ? sub_173898[30:10] : sel_173850[20:0];
  assign shifting_bit_mask__126 = 32'h0000_4000;
  assign sel_173929 = ule_173899 ? sub_173901[30:10] : sel_173853[20:0];
  assign temp__10 = {7'h01, sel_173903, 16'h0000} | shifting_bit_mask__9;
  assign result_sign__864 = 1'h0;
  assign temp__35 = {7'h01, sel_173907, 16'h0000} | shifting_bit_mask__124;
  assign result_sign__865 = 1'h0;
  assign temp__60 = {7'h01, sel_173911, 16'h0000} | shifting_bit_mask__125;
  assign result_sign__866 = 1'h0;
  assign temp__85 = {7'h01, sel_173915, 16'h0000} | shifting_bit_mask__126;
  assign result_sign__867 = 1'h0;
  assign concat_173947 = {sel_173903, result_sign__864};
  assign concat_173952 = {sel_173907, result_sign__865};
  assign concat_173957 = {sel_173911, result_sign__866};
  assign concat_173962 = {sel_173915, result_sign__867};
  assign ule_173966 = temp__10[31:11] <= sel_173920;
  assign sub_173968 = {sel_173920[19:0], 11'h000} - temp__10[30:0];
  assign ule_173969 = temp__35[31:11] <= sel_173923;
  assign sub_173971 = {sel_173923[19:0], 11'h000} - temp__35[30:0];
  assign ule_173972 = temp__60[31:11] <= sel_173926;
  assign sub_173974 = {sel_173926[19:0], 11'h000} - temp__60[30:0];
  assign ule_173975 = temp__85[31:11] <= sel_173929;
  assign sub_173977 = {sel_173929[19:0], 11'h000} - temp__85[30:0];
  assign sel_173979 = ule_173966 ? concat_173947 | 10'h001 : concat_173947;
  assign sel_173983 = ule_173969 ? concat_173952 | 10'h001 : concat_173952;
  assign sel_173987 = ule_173972 ? concat_173957 | 10'h001 : concat_173957;
  assign sel_173991 = ule_173975 ? concat_173962 | 10'h001 : concat_173962;
  assign shifting_bit_mask__10 = 32'h0000_2000;
  assign sel_173996 = ule_173966 ? sub_173968[30:11] : sel_173920[19:0];
  assign shifting_bit_mask__127 = 32'h0000_2000;
  assign sel_173999 = ule_173969 ? sub_173971[30:11] : sel_173923[19:0];
  assign shifting_bit_mask__128 = 32'h0000_2000;
  assign sel_174002 = ule_173972 ? sub_173974[30:11] : sel_173926[19:0];
  assign shifting_bit_mask__129 = 32'h0000_2000;
  assign sel_174005 = ule_173975 ? sub_173977[30:11] : sel_173929[19:0];
  assign temp__11 = {7'h01, sel_173979, 15'h0000} | shifting_bit_mask__10;
  assign result_sign__868 = 1'h0;
  assign temp__36 = {7'h01, sel_173983, 15'h0000} | shifting_bit_mask__127;
  assign result_sign__869 = 1'h0;
  assign temp__61 = {7'h01, sel_173987, 15'h0000} | shifting_bit_mask__128;
  assign result_sign__870 = 1'h0;
  assign temp__86 = {7'h01, sel_173991, 15'h0000} | shifting_bit_mask__129;
  assign result_sign__871 = 1'h0;
  assign concat_174023 = {sel_173979, result_sign__868};
  assign concat_174028 = {sel_173983, result_sign__869};
  assign concat_174033 = {sel_173987, result_sign__870};
  assign concat_174038 = {sel_173991, result_sign__871};
  assign ule_174042 = temp__11[31:12] <= sel_173996;
  assign sub_174044 = {sel_173996[18:0], 12'h000} - temp__11[30:0];
  assign ule_174045 = temp__36[31:12] <= sel_173999;
  assign sub_174047 = {sel_173999[18:0], 12'h000} - temp__36[30:0];
  assign ule_174048 = temp__61[31:12] <= sel_174002;
  assign sub_174050 = {sel_174002[18:0], 12'h000} - temp__61[30:0];
  assign ule_174051 = temp__86[31:12] <= sel_174005;
  assign sub_174053 = {sel_174005[18:0], 12'h000} - temp__86[30:0];
  assign sel_174055 = ule_174042 ? concat_174023 | 11'h001 : concat_174023;
  assign sel_174059 = ule_174045 ? concat_174028 | 11'h001 : concat_174028;
  assign sel_174063 = ule_174048 ? concat_174033 | 11'h001 : concat_174033;
  assign sel_174067 = ule_174051 ? concat_174038 | 11'h001 : concat_174038;
  assign shifting_bit_mask__11 = 32'h0000_1000;
  assign sel_174072 = ule_174042 ? sub_174044[30:12] : sel_173996[18:0];
  assign shifting_bit_mask__130 = 32'h0000_1000;
  assign sel_174075 = ule_174045 ? sub_174047[30:12] : sel_173999[18:0];
  assign shifting_bit_mask__131 = 32'h0000_1000;
  assign sel_174078 = ule_174048 ? sub_174050[30:12] : sel_174002[18:0];
  assign shifting_bit_mask__132 = 32'h0000_1000;
  assign sel_174081 = ule_174051 ? sub_174053[30:12] : sel_174005[18:0];
  assign temp__12 = {7'h01, sel_174055, 14'h0000} | shifting_bit_mask__11;
  assign result_sign__792 = 1'h0;
  assign result_sign__872 = 1'h0;
  assign temp__37 = {7'h01, sel_174059, 14'h0000} | shifting_bit_mask__130;
  assign result_sign__793 = 1'h0;
  assign result_sign__873 = 1'h0;
  assign temp__62 = {7'h01, sel_174063, 14'h0000} | shifting_bit_mask__131;
  assign result_sign__794 = 1'h0;
  assign result_sign__874 = 1'h0;
  assign temp__87 = {7'h01, sel_174067, 14'h0000} | shifting_bit_mask__132;
  assign result_sign__795 = 1'h0;
  assign result_sign__875 = 1'h0;
  assign concat_174104 = {sel_174055, result_sign__872};
  assign concat_174110 = {sel_174059, result_sign__873};
  assign concat_174116 = {sel_174063, result_sign__874};
  assign concat_174122 = {sel_174067, result_sign__875};
  assign ule_174126 = temp__12[31:12] <= {sel_174072, result_sign__792};
  assign result_sign__876 = 1'h0;
  assign sub_174129 = {sel_174072[17:0], 13'h0000} - temp__12[30:0];
  assign ule_174130 = temp__37[31:12] <= {sel_174075, result_sign__793};
  assign result_sign__877 = 1'h0;
  assign sub_174133 = {sel_174075[17:0], 13'h0000} - temp__37[30:0];
  assign ule_174134 = temp__62[31:12] <= {sel_174078, result_sign__794};
  assign result_sign__878 = 1'h0;
  assign sub_174137 = {sel_174078[17:0], 13'h0000} - temp__62[30:0];
  assign ule_174138 = temp__87[31:12] <= {sel_174081, result_sign__795};
  assign result_sign__879 = 1'h0;
  assign sub_174141 = {sel_174081[17:0], 13'h0000} - temp__87[30:0];
  assign sel_174143 = ule_174126 ? concat_174104 | 12'h001 : concat_174104;
  assign sel_174148 = ule_174130 ? concat_174110 | 12'h001 : concat_174110;
  assign sel_174153 = ule_174134 ? concat_174116 | 12'h001 : concat_174116;
  assign sel_174158 = ule_174138 ? concat_174122 | 12'h001 : concat_174122;
  assign shifting_bit_mask__12 = 32'h0000_0800;
  assign sel_174164 = ule_174126 ? sub_174129[30:12] : {sel_174072[17:0], result_sign__876};
  assign shifting_bit_mask__133 = 32'h0000_0800;
  assign sel_174167 = ule_174130 ? sub_174133[30:12] : {sel_174075[17:0], result_sign__877};
  assign shifting_bit_mask__134 = 32'h0000_0800;
  assign sel_174170 = ule_174134 ? sub_174137[30:12] : {sel_174078[17:0], result_sign__878};
  assign shifting_bit_mask__135 = 32'h0000_0800;
  assign sel_174173 = ule_174138 ? sub_174141[30:12] : {sel_174081[17:0], result_sign__879};
  assign temp__13 = {7'h01, sel_174143, 13'h0000} | shifting_bit_mask__12;
  assign result_sign__880 = 1'h0;
  assign temp__38 = {7'h01, sel_174148, 13'h0000} | shifting_bit_mask__133;
  assign result_sign__881 = 1'h0;
  assign temp__63 = {7'h01, sel_174153, 13'h0000} | shifting_bit_mask__134;
  assign result_sign__882 = 1'h0;
  assign temp__88 = {7'h01, sel_174158, 13'h0000} | shifting_bit_mask__135;
  assign result_sign__883 = 1'h0;
  assign concat_174196 = {sel_174143, result_sign__880};
  assign concat_174202 = {sel_174148, result_sign__881};
  assign concat_174208 = {sel_174153, result_sign__882};
  assign concat_174214 = {sel_174158, result_sign__883};
  assign ule_174218 = temp__13[31:11] <= {sel_174164, 2'h0};
  assign sub_174221 = {sel_174164[17:0], 13'h0000} - temp__13[30:0];
  assign ule_174222 = temp__38[31:11] <= {sel_174167, 2'h0};
  assign sub_174225 = {sel_174167[17:0], 13'h0000} - temp__38[30:0];
  assign ule_174226 = temp__63[31:11] <= {sel_174170, 2'h0};
  assign sub_174229 = {sel_174170[17:0], 13'h0000} - temp__63[30:0];
  assign ule_174230 = temp__88[31:11] <= {sel_174173, 2'h0};
  assign sub_174233 = {sel_174173[17:0], 13'h0000} - temp__88[30:0];
  assign sel_174235 = ule_174218 ? concat_174196 | 13'h0001 : concat_174196;
  assign sel_174240 = ule_174222 ? concat_174202 | 13'h0001 : concat_174202;
  assign sel_174245 = ule_174226 ? concat_174208 | 13'h0001 : concat_174208;
  assign sel_174250 = ule_174230 ? concat_174214 | 13'h0001 : concat_174214;
  assign shifting_bit_mask__13 = 32'h0000_0400;
  assign sel_174256 = ule_174218 ? sub_174221[30:11] : {sel_174164[17:0], 2'h0};
  assign shifting_bit_mask__136 = 32'h0000_0400;
  assign sel_174259 = ule_174222 ? sub_174225[30:11] : {sel_174167[17:0], 2'h0};
  assign shifting_bit_mask__137 = 32'h0000_0400;
  assign sel_174262 = ule_174226 ? sub_174229[30:11] : {sel_174170[17:0], 2'h0};
  assign shifting_bit_mask__138 = 32'h0000_0400;
  assign sel_174265 = ule_174230 ? sub_174233[30:11] : {sel_174173[17:0], 2'h0};
  assign temp__14 = {7'h01, sel_174235, 12'h000} | shifting_bit_mask__13;
  assign result_sign__884 = 1'h0;
  assign temp__39 = {7'h01, sel_174240, 12'h000} | shifting_bit_mask__136;
  assign result_sign__885 = 1'h0;
  assign temp__64 = {7'h01, sel_174245, 12'h000} | shifting_bit_mask__137;
  assign result_sign__886 = 1'h0;
  assign temp__89 = {7'h01, sel_174250, 12'h000} | shifting_bit_mask__138;
  assign result_sign__887 = 1'h0;
  assign concat_174288 = {sel_174235, result_sign__884};
  assign concat_174294 = {sel_174240, result_sign__885};
  assign concat_174300 = {sel_174245, result_sign__886};
  assign concat_174306 = {sel_174250, result_sign__887};
  assign ule_174310 = temp__14[31:10] <= {sel_174256, 2'h0};
  assign sub_174313 = {sel_174256[18:0], 12'h000} - temp__14[30:0];
  assign ule_174314 = temp__39[31:10] <= {sel_174259, 2'h0};
  assign sub_174317 = {sel_174259[18:0], 12'h000} - temp__39[30:0];
  assign ule_174318 = temp__64[31:10] <= {sel_174262, 2'h0};
  assign sub_174321 = {sel_174262[18:0], 12'h000} - temp__64[30:0];
  assign ule_174322 = temp__89[31:10] <= {sel_174265, 2'h0};
  assign sub_174325 = {sel_174265[18:0], 12'h000} - temp__89[30:0];
  assign sel_174327 = ule_174310 ? concat_174288 | 14'h0001 : concat_174288;
  assign sel_174332 = ule_174314 ? concat_174294 | 14'h0001 : concat_174294;
  assign sel_174337 = ule_174318 ? concat_174300 | 14'h0001 : concat_174300;
  assign sel_174342 = ule_174322 ? concat_174306 | 14'h0001 : concat_174306;
  assign shifting_bit_mask__14 = 32'h0000_0200;
  assign sel_174348 = ule_174310 ? sub_174313[30:10] : {sel_174256[18:0], 2'h0};
  assign shifting_bit_mask__139 = 32'h0000_0200;
  assign sel_174351 = ule_174314 ? sub_174317[30:10] : {sel_174259[18:0], 2'h0};
  assign shifting_bit_mask__140 = 32'h0000_0200;
  assign sel_174354 = ule_174318 ? sub_174321[30:10] : {sel_174262[18:0], 2'h0};
  assign shifting_bit_mask__141 = 32'h0000_0200;
  assign sel_174357 = ule_174322 ? sub_174325[30:10] : {sel_174265[18:0], 2'h0};
  assign temp__15 = {7'h01, sel_174327, 11'h000} | shifting_bit_mask__14;
  assign result_sign__888 = 1'h0;
  assign temp__40 = {7'h01, sel_174332, 11'h000} | shifting_bit_mask__139;
  assign result_sign__889 = 1'h0;
  assign temp__65 = {7'h01, sel_174337, 11'h000} | shifting_bit_mask__140;
  assign result_sign__890 = 1'h0;
  assign temp__90 = {7'h01, sel_174342, 11'h000} | shifting_bit_mask__141;
  assign result_sign__891 = 1'h0;
  assign concat_174380 = {sel_174327, result_sign__888};
  assign concat_174386 = {sel_174332, result_sign__889};
  assign concat_174392 = {sel_174337, result_sign__890};
  assign concat_174398 = {sel_174342, result_sign__891};
  assign ule_174402 = temp__15[31:9] <= {sel_174348, 2'h0};
  assign sub_174405 = {sel_174348[19:0], 11'h000} - temp__15[30:0];
  assign ule_174406 = temp__40[31:9] <= {sel_174351, 2'h0};
  assign sub_174409 = {sel_174351[19:0], 11'h000} - temp__40[30:0];
  assign ule_174410 = temp__65[31:9] <= {sel_174354, 2'h0};
  assign sub_174413 = {sel_174354[19:0], 11'h000} - temp__65[30:0];
  assign ule_174414 = temp__90[31:9] <= {sel_174357, 2'h0};
  assign sub_174417 = {sel_174357[19:0], 11'h000} - temp__90[30:0];
  assign sel_174419 = ule_174402 ? concat_174380 | 15'h0001 : concat_174380;
  assign sel_174424 = ule_174406 ? concat_174386 | 15'h0001 : concat_174386;
  assign sel_174429 = ule_174410 ? concat_174392 | 15'h0001 : concat_174392;
  assign sel_174434 = ule_174414 ? concat_174398 | 15'h0001 : concat_174398;
  assign shifting_bit_mask__15 = 32'h0000_0100;
  assign sel_174440 = ule_174402 ? sub_174405[30:9] : {sel_174348[19:0], 2'h0};
  assign shifting_bit_mask__142 = 32'h0000_0100;
  assign sel_174443 = ule_174406 ? sub_174409[30:9] : {sel_174351[19:0], 2'h0};
  assign shifting_bit_mask__143 = 32'h0000_0100;
  assign sel_174446 = ule_174410 ? sub_174413[30:9] : {sel_174354[19:0], 2'h0};
  assign shifting_bit_mask__144 = 32'h0000_0100;
  assign sel_174449 = ule_174414 ? sub_174417[30:9] : {sel_174357[19:0], 2'h0};
  assign temp__16 = {7'h01, sel_174419, 10'h000} | shifting_bit_mask__15;
  assign result_sign__892 = 1'h0;
  assign temp__41 = {7'h01, sel_174424, 10'h000} | shifting_bit_mask__142;
  assign result_sign__893 = 1'h0;
  assign temp__66 = {7'h01, sel_174429, 10'h000} | shifting_bit_mask__143;
  assign result_sign__894 = 1'h0;
  assign temp__91 = {7'h01, sel_174434, 10'h000} | shifting_bit_mask__144;
  assign result_sign__895 = 1'h0;
  assign concat_174472 = {sel_174419, result_sign__892};
  assign concat_174478 = {sel_174424, result_sign__893};
  assign concat_174484 = {sel_174429, result_sign__894};
  assign concat_174490 = {sel_174434, result_sign__895};
  assign ule_174494 = temp__16[31:8] <= {sel_174440, 2'h0};
  assign sub_174497 = {sel_174440[20:0], 10'h000} - temp__16[30:0];
  assign ule_174498 = temp__41[31:8] <= {sel_174443, 2'h0};
  assign sub_174501 = {sel_174443[20:0], 10'h000} - temp__41[30:0];
  assign ule_174502 = temp__66[31:8] <= {sel_174446, 2'h0};
  assign sub_174505 = {sel_174446[20:0], 10'h000} - temp__66[30:0];
  assign ule_174506 = temp__91[31:8] <= {sel_174449, 2'h0};
  assign sub_174509 = {sel_174449[20:0], 10'h000} - temp__91[30:0];
  assign sel_174511 = ule_174494 ? concat_174472 | 16'h0001 : concat_174472;
  assign sel_174516 = ule_174498 ? concat_174478 | 16'h0001 : concat_174478;
  assign sel_174521 = ule_174502 ? concat_174484 | 16'h0001 : concat_174484;
  assign sel_174526 = ule_174506 ? concat_174490 | 16'h0001 : concat_174490;
  assign shifting_bit_mask__16 = 32'h0000_0080;
  assign sel_174532 = ule_174494 ? sub_174497[30:8] : {sel_174440[20:0], 2'h0};
  assign shifting_bit_mask__145 = 32'h0000_0080;
  assign sel_174535 = ule_174498 ? sub_174501[30:8] : {sel_174443[20:0], 2'h0};
  assign shifting_bit_mask__146 = 32'h0000_0080;
  assign sel_174538 = ule_174502 ? sub_174505[30:8] : {sel_174446[20:0], 2'h0};
  assign shifting_bit_mask__147 = 32'h0000_0080;
  assign sel_174541 = ule_174506 ? sub_174509[30:8] : {sel_174449[20:0], 2'h0};
  assign temp__17 = {7'h01, sel_174511, 9'h000} | shifting_bit_mask__16;
  assign result_sign__896 = 1'h0;
  assign temp__42 = {7'h01, sel_174516, 9'h000} | shifting_bit_mask__145;
  assign result_sign__897 = 1'h0;
  assign temp__67 = {7'h01, sel_174521, 9'h000} | shifting_bit_mask__146;
  assign result_sign__898 = 1'h0;
  assign temp__92 = {7'h01, sel_174526, 9'h000} | shifting_bit_mask__147;
  assign result_sign__899 = 1'h0;
  assign concat_174564 = {sel_174511, result_sign__896};
  assign concat_174570 = {sel_174516, result_sign__897};
  assign concat_174576 = {sel_174521, result_sign__898};
  assign concat_174582 = {sel_174526, result_sign__899};
  assign ule_174586 = temp__17[31:7] <= {sel_174532, 2'h0};
  assign sub_174589 = {sel_174532[21:0], 9'h000} - temp__17[30:0];
  assign ule_174590 = temp__42[31:7] <= {sel_174535, 2'h0};
  assign sub_174593 = {sel_174535[21:0], 9'h000} - temp__42[30:0];
  assign ule_174594 = temp__67[31:7] <= {sel_174538, 2'h0};
  assign sub_174597 = {sel_174538[21:0], 9'h000} - temp__67[30:0];
  assign ule_174598 = temp__92[31:7] <= {sel_174541, 2'h0};
  assign sub_174601 = {sel_174541[21:0], 9'h000} - temp__92[30:0];
  assign sel_174603 = ule_174586 ? concat_174564 | 17'h0_0001 : concat_174564;
  assign x_bexp__652 = 8'h00;
  assign sel_174608 = ule_174590 ? concat_174570 | 17'h0_0001 : concat_174570;
  assign x_bexp__653 = 8'h00;
  assign sel_174613 = ule_174594 ? concat_174576 | 17'h0_0001 : concat_174576;
  assign x_bexp__654 = 8'h00;
  assign sel_174618 = ule_174598 ? concat_174582 | 17'h0_0001 : concat_174582;
  assign x_bexp__655 = 8'h00;
  assign shifting_bit_mask__17 = 32'h0000_0040;
  assign sel_174624 = ule_174586 ? sub_174589[30:7] : {sel_174532[21:0], 2'h0};
  assign shifting_bit_mask__148 = 32'h0000_0040;
  assign sel_174627 = ule_174590 ? sub_174593[30:7] : {sel_174535[21:0], 2'h0};
  assign shifting_bit_mask__149 = 32'h0000_0040;
  assign sel_174630 = ule_174594 ? sub_174597[30:7] : {sel_174538[21:0], 2'h0};
  assign shifting_bit_mask__150 = 32'h0000_0040;
  assign sel_174633 = ule_174598 ? sub_174601[30:7] : {sel_174541[21:0], 2'h0};
  assign temp__18 = {7'h01, sel_174603, x_bexp__652} | shifting_bit_mask__17;
  assign result_sign__900 = 1'h0;
  assign x_bexp__657 = 8'h00;
  assign temp__43 = {7'h01, sel_174608, x_bexp__653} | shifting_bit_mask__148;
  assign result_sign__901 = 1'h0;
  assign x_bexp__659 = 8'h00;
  assign temp__68 = {7'h01, sel_174613, x_bexp__654} | shifting_bit_mask__149;
  assign result_sign__902 = 1'h0;
  assign x_bexp__661 = 8'h00;
  assign temp__93 = {7'h01, sel_174618, x_bexp__655} | shifting_bit_mask__150;
  assign result_sign__903 = 1'h0;
  assign x_bexp__663 = 8'h00;
  assign concat_174656 = {sel_174603, result_sign__900};
  assign concat_174662 = {sel_174608, result_sign__901};
  assign concat_174668 = {sel_174613, result_sign__902};
  assign concat_174674 = {sel_174618, result_sign__903};
  assign ule_174678 = temp__18[31:6] <= {sel_174624, 2'h0};
  assign sub_174681 = {sel_174624[22:0], x_bexp__657} - temp__18[30:0];
  assign ule_174682 = temp__43[31:6] <= {sel_174627, 2'h0};
  assign sub_174685 = {sel_174627[22:0], x_bexp__659} - temp__43[30:0];
  assign ule_174686 = temp__68[31:6] <= {sel_174630, 2'h0};
  assign sub_174689 = {sel_174630[22:0], x_bexp__661} - temp__68[30:0];
  assign ule_174690 = temp__93[31:6] <= {sel_174633, 2'h0};
  assign sub_174693 = {sel_174633[22:0], x_bexp__663} - temp__93[30:0];
  assign sel_174695 = ule_174678 ? concat_174656 | 18'h0_0001 : concat_174656;
  assign sel_174700 = ule_174682 ? concat_174662 | 18'h0_0001 : concat_174662;
  assign sel_174705 = ule_174686 ? concat_174668 | 18'h0_0001 : concat_174668;
  assign sel_174710 = ule_174690 ? concat_174674 | 18'h0_0001 : concat_174674;
  assign shifting_bit_mask__18 = 32'h0000_0020;
  assign sel_174716 = ule_174678 ? sub_174681[30:6] : {sel_174624[22:0], 2'h0};
  assign shifting_bit_mask__151 = 32'h0000_0020;
  assign sel_174719 = ule_174682 ? sub_174685[30:6] : {sel_174627[22:0], 2'h0};
  assign shifting_bit_mask__152 = 32'h0000_0020;
  assign sel_174722 = ule_174686 ? sub_174689[30:6] : {sel_174630[22:0], 2'h0};
  assign shifting_bit_mask__153 = 32'h0000_0020;
  assign sel_174725 = ule_174690 ? sub_174693[30:6] : {sel_174633[22:0], 2'h0};
  assign temp__19 = {7'h01, sel_174695, 7'h00} | shifting_bit_mask__18;
  assign result_sign__904 = 1'h0;
  assign temp__44 = {7'h01, sel_174700, 7'h00} | shifting_bit_mask__151;
  assign result_sign__905 = 1'h0;
  assign temp__69 = {7'h01, sel_174705, 7'h00} | shifting_bit_mask__152;
  assign result_sign__906 = 1'h0;
  assign temp__94 = {7'h01, sel_174710, 7'h00} | shifting_bit_mask__153;
  assign result_sign__907 = 1'h0;
  assign concat_174748 = {sel_174695, result_sign__904};
  assign concat_174754 = {sel_174700, result_sign__905};
  assign concat_174760 = {sel_174705, result_sign__906};
  assign concat_174766 = {sel_174710, result_sign__907};
  assign ule_174770 = temp__19[31:5] <= {sel_174716, 2'h0};
  assign sub_174773 = {sel_174716[23:0], 7'h00} - temp__19[30:0];
  assign ule_174774 = temp__44[31:5] <= {sel_174719, 2'h0};
  assign sub_174777 = {sel_174719[23:0], 7'h00} - temp__44[30:0];
  assign ule_174778 = temp__69[31:5] <= {sel_174722, 2'h0};
  assign sub_174781 = {sel_174722[23:0], 7'h00} - temp__69[30:0];
  assign ule_174782 = temp__94[31:5] <= {sel_174725, 2'h0};
  assign sub_174785 = {sel_174725[23:0], 7'h00} - temp__94[30:0];
  assign sel_174787 = ule_174770 ? concat_174748 | 19'h0_0001 : concat_174748;
  assign sel_174792 = ule_174774 ? concat_174754 | 19'h0_0001 : concat_174754;
  assign sel_174797 = ule_174778 ? concat_174760 | 19'h0_0001 : concat_174760;
  assign sel_174802 = ule_174782 ? concat_174766 | 19'h0_0001 : concat_174766;
  assign shifting_bit_mask__19 = 32'h0000_0010;
  assign sel_174808 = ule_174770 ? sub_174773[30:5] : {sel_174716[23:0], 2'h0};
  assign shifting_bit_mask__154 = 32'h0000_0010;
  assign sel_174811 = ule_174774 ? sub_174777[30:5] : {sel_174719[23:0], 2'h0};
  assign shifting_bit_mask__155 = 32'h0000_0010;
  assign sel_174814 = ule_174778 ? sub_174781[30:5] : {sel_174722[23:0], 2'h0};
  assign shifting_bit_mask__156 = 32'h0000_0010;
  assign sel_174817 = ule_174782 ? sub_174785[30:5] : {sel_174725[23:0], 2'h0};
  assign temp__20 = {7'h01, sel_174787, 6'h00} | shifting_bit_mask__19;
  assign result_sign__908 = 1'h0;
  assign temp__45 = {7'h01, sel_174792, 6'h00} | shifting_bit_mask__154;
  assign result_sign__909 = 1'h0;
  assign temp__70 = {7'h01, sel_174797, 6'h00} | shifting_bit_mask__155;
  assign result_sign__910 = 1'h0;
  assign temp__95 = {7'h01, sel_174802, 6'h00} | shifting_bit_mask__156;
  assign result_sign__911 = 1'h0;
  assign concat_174840 = {sel_174787, result_sign__908};
  assign concat_174846 = {sel_174792, result_sign__909};
  assign concat_174852 = {sel_174797, result_sign__910};
  assign concat_174858 = {sel_174802, result_sign__911};
  assign ule_174862 = temp__20[31:4] <= {sel_174808, 2'h0};
  assign sub_174865 = {sel_174808[24:0], 6'h00} - temp__20[30:0];
  assign ule_174866 = temp__45[31:4] <= {sel_174811, 2'h0};
  assign sub_174869 = {sel_174811[24:0], 6'h00} - temp__45[30:0];
  assign ule_174870 = temp__70[31:4] <= {sel_174814, 2'h0};
  assign sub_174873 = {sel_174814[24:0], 6'h00} - temp__70[30:0];
  assign ule_174874 = temp__95[31:4] <= {sel_174817, 2'h0};
  assign sub_174877 = {sel_174817[24:0], 6'h00} - temp__95[30:0];
  assign sel_174879 = ule_174862 ? concat_174840 | 20'h0_0001 : concat_174840;
  assign sel_174884 = ule_174866 ? concat_174846 | 20'h0_0001 : concat_174846;
  assign sel_174889 = ule_174870 ? concat_174852 | 20'h0_0001 : concat_174852;
  assign sel_174894 = ule_174874 ? concat_174858 | 20'h0_0001 : concat_174858;
  assign shifting_bit_mask__20 = 32'h0000_0008;
  assign sel_174900 = ule_174862 ? sub_174865[30:4] : {sel_174808[24:0], 2'h0};
  assign shifting_bit_mask__157 = 32'h0000_0008;
  assign sel_174903 = ule_174866 ? sub_174869[30:4] : {sel_174811[24:0], 2'h0};
  assign shifting_bit_mask__158 = 32'h0000_0008;
  assign sel_174906 = ule_174870 ? sub_174873[30:4] : {sel_174814[24:0], 2'h0};
  assign shifting_bit_mask__159 = 32'h0000_0008;
  assign sel_174909 = ule_174874 ? sub_174877[30:4] : {sel_174817[24:0], 2'h0};
  assign temp__21 = {7'h01, sel_174879, 5'h00} | shifting_bit_mask__20;
  assign result_sign__912 = 1'h0;
  assign temp__46 = {7'h01, sel_174884, 5'h00} | shifting_bit_mask__157;
  assign result_sign__913 = 1'h0;
  assign temp__71 = {7'h01, sel_174889, 5'h00} | shifting_bit_mask__158;
  assign result_sign__914 = 1'h0;
  assign temp__96 = {7'h01, sel_174894, 5'h00} | shifting_bit_mask__159;
  assign result_sign__915 = 1'h0;
  assign concat_174932 = {sel_174879, result_sign__912};
  assign concat_174938 = {sel_174884, result_sign__913};
  assign concat_174944 = {sel_174889, result_sign__914};
  assign concat_174950 = {sel_174894, result_sign__915};
  assign ule_174954 = temp__21[31:3] <= {sel_174900, 2'h0};
  assign sub_174957 = {sel_174900[25:0], 5'h00} - temp__21[30:0];
  assign ule_174958 = temp__46[31:3] <= {sel_174903, 2'h0};
  assign sub_174961 = {sel_174903[25:0], 5'h00} - temp__46[30:0];
  assign ule_174962 = temp__71[31:3] <= {sel_174906, 2'h0};
  assign sub_174965 = {sel_174906[25:0], 5'h00} - temp__71[30:0];
  assign ule_174966 = temp__96[31:3] <= {sel_174909, 2'h0};
  assign sub_174969 = {sel_174909[25:0], 5'h00} - temp__96[30:0];
  assign sel_174971 = ule_174954 ? concat_174932 | 21'h00_0001 : concat_174932;
  assign sel_174976 = ule_174958 ? concat_174938 | 21'h00_0001 : concat_174938;
  assign sel_174981 = ule_174962 ? concat_174944 | 21'h00_0001 : concat_174944;
  assign sel_174986 = ule_174966 ? concat_174950 | 21'h00_0001 : concat_174950;
  assign shifting_bit_mask__21 = 32'h0000_0004;
  assign sel_174992 = ule_174954 ? sub_174957[30:3] : {sel_174900[25:0], 2'h0};
  assign shifting_bit_mask__160 = 32'h0000_0004;
  assign sel_174995 = ule_174958 ? sub_174961[30:3] : {sel_174903[25:0], 2'h0};
  assign shifting_bit_mask__161 = 32'h0000_0004;
  assign sel_174998 = ule_174962 ? sub_174965[30:3] : {sel_174906[25:0], 2'h0};
  assign shifting_bit_mask__162 = 32'h0000_0004;
  assign sel_175001 = ule_174966 ? sub_174969[30:3] : {sel_174909[25:0], 2'h0};
  assign temp__22 = {7'h01, sel_174971, 4'h0} | shifting_bit_mask__21;
  assign result_sign__916 = 1'h0;
  assign temp__47 = {7'h01, sel_174976, 4'h0} | shifting_bit_mask__160;
  assign result_sign__917 = 1'h0;
  assign temp__72 = {7'h01, sel_174981, 4'h0} | shifting_bit_mask__161;
  assign result_sign__918 = 1'h0;
  assign temp__97 = {7'h01, sel_174986, 4'h0} | shifting_bit_mask__162;
  assign result_sign__919 = 1'h0;
  assign concat_175024 = {sel_174971, result_sign__916};
  assign concat_175030 = {sel_174976, result_sign__917};
  assign concat_175036 = {sel_174981, result_sign__918};
  assign concat_175042 = {sel_174986, result_sign__919};
  assign ule_175046 = temp__22[31:2] <= {sel_174992, 2'h0};
  assign sub_175049 = {sel_174992[26:0], 4'h0} - temp__22[30:0];
  assign ule_175050 = temp__47[31:2] <= {sel_174995, 2'h0};
  assign sub_175053 = {sel_174995[26:0], 4'h0} - temp__47[30:0];
  assign ule_175054 = temp__72[31:2] <= {sel_174998, 2'h0};
  assign sub_175057 = {sel_174998[26:0], 4'h0} - temp__72[30:0];
  assign ule_175058 = temp__97[31:2] <= {sel_175001, 2'h0};
  assign sub_175061 = {sel_175001[26:0], 4'h0} - temp__97[30:0];
  assign sel_175063 = ule_175046 ? concat_175024 | 22'h00_0001 : concat_175024;
  assign sel_175068 = ule_175050 ? concat_175030 | 22'h00_0001 : concat_175030;
  assign sel_175073 = ule_175054 ? concat_175036 | 22'h00_0001 : concat_175036;
  assign sel_175078 = ule_175058 ? concat_175042 | 22'h00_0001 : concat_175042;
  assign shifting_bit_mask__22 = 32'h0000_0002;
  assign sel_175084 = ule_175046 ? sub_175049[30:2] : {sel_174992[26:0], 2'h0};
  assign shifting_bit_mask__163 = 32'h0000_0002;
  assign sel_175087 = ule_175050 ? sub_175053[30:2] : {sel_174995[26:0], 2'h0};
  assign shifting_bit_mask__164 = 32'h0000_0002;
  assign sel_175090 = ule_175054 ? sub_175057[30:2] : {sel_174998[26:0], 2'h0};
  assign shifting_bit_mask__165 = 32'h0000_0002;
  assign sel_175093 = ule_175058 ? sub_175061[30:2] : {sel_175001[26:0], 2'h0};
  assign temp__23 = {7'h01, sel_175063, 3'h0} | shifting_bit_mask__22;
  assign result_sign__920 = 1'h0;
  assign temp__48 = {7'h01, sel_175068, 3'h0} | shifting_bit_mask__163;
  assign result_sign__921 = 1'h0;
  assign temp__73 = {7'h01, sel_175073, 3'h0} | shifting_bit_mask__164;
  assign result_sign__922 = 1'h0;
  assign temp__98 = {7'h01, sel_175078, 3'h0} | shifting_bit_mask__165;
  assign result_sign__923 = 1'h0;
  assign scaled_fixed_point_x__50 = {sel_175084, 2'h0};
  assign concat_175116 = {sel_175063, result_sign__920};
  assign scaled_fixed_point_x__101 = {sel_175087, 2'h0};
  assign concat_175122 = {sel_175068, result_sign__921};
  assign scaled_fixed_point_x__155 = {sel_175090, 2'h0};
  assign concat_175128 = {sel_175073, result_sign__922};
  assign scaled_fixed_point_x__209 = {sel_175093, 2'h0};
  assign concat_175134 = {sel_175078, result_sign__923};
  assign ule_175138 = temp__23[31:1] <= scaled_fixed_point_x__50;
  assign sub_175141 = {sel_175084[27:0], 3'h0} - temp__23[30:0];
  assign ule_175142 = temp__48[31:1] <= scaled_fixed_point_x__101;
  assign sub_175145 = {sel_175087[27:0], 3'h0} - temp__48[30:0];
  assign ule_175146 = temp__73[31:1] <= scaled_fixed_point_x__155;
  assign sub_175149 = {sel_175090[27:0], 3'h0} - temp__73[30:0];
  assign ule_175150 = temp__98[31:1] <= scaled_fixed_point_x__209;
  assign sub_175153 = {sel_175093[27:0], 3'h0} - temp__98[30:0];
  assign sel_175155 = ule_175138 ? concat_175116 | 23'h00_0001 : concat_175116;
  assign sel_175160 = ule_175142 ? concat_175122 | 23'h00_0001 : concat_175122;
  assign sel_175165 = ule_175146 ? concat_175128 | 23'h00_0001 : concat_175128;
  assign sel_175170 = ule_175150 ? concat_175134 | 23'h00_0001 : concat_175134;
  assign shifting_bit_mask__23 = 32'h0000_0001;
  assign sel_175176 = ule_175138 ? sub_175141[30:1] : {sel_175084[27:0], 2'h0};
  assign result_sign__924 = 1'h0;
  assign shifting_bit_mask__166 = 32'h0000_0001;
  assign sel_175181 = ule_175142 ? sub_175145[30:1] : {sel_175087[27:0], 2'h0};
  assign result_sign__925 = 1'h0;
  assign shifting_bit_mask__167 = 32'h0000_0001;
  assign sel_175186 = ule_175146 ? sub_175149[30:1] : {sel_175090[27:0], 2'h0};
  assign result_sign__926 = 1'h0;
  assign shifting_bit_mask__168 = 32'h0000_0001;
  assign sel_175191 = ule_175150 ? sub_175153[30:1] : {sel_175093[27:0], 2'h0};
  assign result_sign__927 = 1'h0;
  assign temp__24 = {7'h01, sel_175155, 2'h0} | shifting_bit_mask__23;
  assign scaled_fixed_point_x__53 = {sel_175176, 2'h0};
  assign concat_175196 = {sel_175155, result_sign__924};
  assign temp__49 = {7'h01, sel_175160, 2'h0} | shifting_bit_mask__166;
  assign scaled_fixed_point_x__104 = {sel_175181, 2'h0};
  assign concat_175200 = {sel_175160, result_sign__925};
  assign temp__74 = {7'h01, sel_175165, 2'h0} | shifting_bit_mask__167;
  assign scaled_fixed_point_x__158 = {sel_175186, 2'h0};
  assign concat_175204 = {sel_175165, result_sign__926};
  assign temp__99 = {7'h01, sel_175170, 2'h0} | shifting_bit_mask__168;
  assign scaled_fixed_point_x__212 = {sel_175191, 2'h0};
  assign concat_175208 = {sel_175170, result_sign__927};
  assign ule_175212 = temp__24 <= scaled_fixed_point_x__53;
  assign ule_175216 = temp__49 <= scaled_fixed_point_x__104;
  assign ule_175220 = temp__74 <= scaled_fixed_point_x__158;
  assign ule_175224 = temp__99 <= scaled_fixed_point_x__212;
  assign concat_175226 = {sel_175176[28:0], 2'h0};
  assign sel_175229 = ule_175212 ? concat_175196 | 24'h00_0001 : concat_175196;
  assign concat_175231 = {sel_175181[28:0], 2'h0};
  assign sel_175234 = ule_175216 ? concat_175200 | 24'h00_0001 : concat_175200;
  assign concat_175236 = {sel_175186[28:0], 2'h0};
  assign sel_175239 = ule_175220 ? concat_175204 | 24'h00_0001 : concat_175204;
  assign concat_175241 = {sel_175191[28:0], 2'h0};
  assign sel_175244 = ule_175224 ? concat_175208 | 24'h00_0001 : concat_175208;
  assign sub_175246 = concat_175226 - temp__24[30:0];
  assign sub_175249 = concat_175231 - temp__49[30:0];
  assign sub_175252 = concat_175236 - temp__74[30:0];
  assign sub_175255 = concat_175241 - temp__99[30:0];
  assign scaled_fixed_point_x__54 = ule_175212 ? sub_175246 : concat_175226;
  assign add_175262 = {2'h1, sel_175229} + {25'h000_0000, ule_175212};
  assign scaled_fixed_point_x__105 = ule_175216 ? sub_175249 : concat_175231;
  assign add_175267 = {2'h1, sel_175234} + {25'h000_0000, ule_175216};
  assign scaled_fixed_point_x__159 = ule_175220 ? sub_175252 : concat_175236;
  assign add_175272 = {2'h1, sel_175239} + {25'h000_0000, ule_175220};
  assign scaled_fixed_point_x__213 = ule_175224 ? sub_175255 : concat_175241;
  assign add_175277 = {2'h1, sel_175244} + {25'h000_0000, ule_175224};
  assign bit_slice_175281 = uexp[7:2];
  assign bit_slice_175285 = uexp__1[7:2];
  assign bit_slice_175289 = uexp__2[7:2];
  assign bit_slice_175293 = uexp__3[7:2];
  assign sel_175294 = scaled_fixed_point_x__54 != 31'h0000_0000 ? add_175262[25:1] : {2'h1, sel_175229[23:1]};
  assign sel_175297 = scaled_fixed_point_x__105 != 31'h0000_0000 ? add_175267[25:1] : {2'h1, sel_175234[23:1]};
  assign sel_175300 = scaled_fixed_point_x__159 != 31'h0000_0000 ? add_175272[25:1] : {2'h1, sel_175239[23:1]};
  assign sel_175303 = scaled_fixed_point_x__213 != 31'h0000_0000 ? add_175277[25:1] : {2'h1, sel_175244[23:1]};
  assign result_sign__1120 = 1'h0;
  assign add_175309 = {{1{bit_slice_175281[5]}}, bit_slice_175281} + 7'h3f;
  assign result_sign__1121 = 1'h0;
  assign add_175314 = {{1{bit_slice_175285[5]}}, bit_slice_175285} + 7'h3f;
  assign result_sign__1122 = 1'h0;
  assign add_175319 = {{1{bit_slice_175289[5]}}, bit_slice_175289} + 7'h3f;
  assign result_sign__1123 = 1'h0;
  assign add_175324 = {{1{bit_slice_175293[5]}}, bit_slice_175293} + 7'h3f;
  assign high_exp__141 = 8'hff;
  assign result_fraction__541 = 23'h00_0000;
  assign high_exp__207 = 8'hff;
  assign result_fraction__608 = 23'h00_0000;
  assign high_exp__275 = 8'hff;
  assign result_fraction__675 = 23'h00_0000;
  assign high_exp__349 = 8'hff;
  assign result_fraction__754 = 23'h00_0000;
  assign eq_175342 = result_exponent__19 == high_exp__141;
  assign eq_175343 = result_fraction__117 == result_fraction__541;
  assign add_175344 = {7'h00, sel_175294[24:23]} + {result_sign__1120, add_175309, uexp[1]};
  assign eq_175345 = result_exponent__38 == high_exp__207;
  assign eq_175346 = result_fraction__234 == result_fraction__608;
  assign add_175347 = {7'h00, sel_175297[24:23]} + {result_sign__1121, add_175314, uexp__1[1]};
  assign eq_175348 = result_exponent__57 == high_exp__275;
  assign eq_175349 = result_fraction__351 == result_fraction__675;
  assign add_175350 = {7'h00, sel_175300[24:23]} + {result_sign__1122, add_175319, uexp__2[1]};
  assign eq_175351 = result_exponent__76 == high_exp__349;
  assign eq_175352 = result_fraction__468 == result_fraction__754;
  assign add_175353 = {7'h00, sel_175303[24:23]} + {result_sign__1123, add_175324, uexp__3[1]};
  assign result_fraction__542 = 23'h00_0000;
  assign result_fraction__609 = 23'h00_0000;
  assign result_fraction__676 = 23'h00_0000;
  assign result_fraction__755 = 23'h00_0000;
  assign and_175368 = eq_175342 & eq_175343;
  assign x_bexp__828 = 8'h00;
  assign and_175374 = eq_175345 & eq_175346;
  assign x_bexp__829 = 8'h00;
  assign and_175380 = eq_175348 & eq_175349;
  assign x_bexp__830 = 8'h00;
  assign and_175386 = eq_175351 & eq_175352;
  assign x_bexp__831 = 8'h00;
  assign and_175390 = eq_175342 & result_fraction__117 != result_fraction__542;
  assign x_bexp__593 = 8'h00;
  assign high_exp__142 = 8'hff;
  assign nan_fraction__106 = 23'h40_0000;
  assign ne_175397 = result_exponent__19 != x_bexp__828;
  assign and_175398 = eq_175345 & result_fraction__234 != result_fraction__609;
  assign x_bexp__611 = 8'h00;
  assign high_exp__208 = 8'hff;
  assign nan_fraction__133 = 23'h40_0000;
  assign ne_175405 = result_exponent__38 != x_bexp__829;
  assign and_175406 = eq_175348 & result_fraction__351 != result_fraction__676;
  assign x_bexp__629 = 8'h00;
  assign high_exp__276 = 8'hff;
  assign nan_fraction__162 = 23'h40_0000;
  assign ne_175413 = result_exponent__57 != x_bexp__830;
  assign and_175414 = eq_175351 & result_fraction__468 != result_fraction__755;
  assign x_bexp__647 = 8'h00;
  assign high_exp__350 = 8'hff;
  assign nan_fraction__191 = 23'h40_0000;
  assign ne_175421 = result_exponent__76 != x_bexp__831;
  assign pixel_val = {ne_175397 & ~(and_175390 | ~(~(eq_175342 & eq_175343) & add_175344[8])), result_exponent__19 == x_bexp__593 ? result_exponent__19 : (and_175390 ? high_exp__142 : (and_175368 ? result_exponent__19 : add_175344[7:0])), (and_175390 ? nan_fraction__106 : (and_175368 ? result_fraction__117 : sel_175294[22:0])) & {23{ne_175397}}};
  assign pixel_val__1 = {ne_175405 & ~(and_175398 | ~(~(eq_175345 & eq_175346) & add_175347[8])), result_exponent__38 == x_bexp__611 ? result_exponent__38 : (and_175398 ? high_exp__208 : (and_175374 ? result_exponent__38 : add_175347[7:0])), (and_175398 ? nan_fraction__133 : (and_175374 ? result_fraction__234 : sel_175297[22:0])) & {23{ne_175405}}};
  assign pixel_val__2 = {ne_175413 & ~(and_175406 | ~(~(eq_175348 & eq_175349) & add_175350[8])), result_exponent__57 == x_bexp__629 ? result_exponent__57 : (and_175406 ? high_exp__276 : (and_175380 ? result_exponent__57 : add_175350[7:0])), (and_175406 ? nan_fraction__162 : (and_175380 ? result_fraction__351 : sel_175300[22:0])) & {23{ne_175413}}};
  assign pixel_val__3 = {ne_175421 & ~(and_175414 | ~(~(eq_175351 & eq_175352) & add_175353[8])), result_exponent__76 == x_bexp__647 ? result_exponent__76 : (and_175414 ? high_exp__350 : (and_175386 ? result_exponent__76 : add_175353[7:0])), (and_175414 ? nan_fraction__191 : (and_175386 ? result_fraction__468 : sel_175303[22:0])) & {23{ne_175421}}};
  assign array_175531[0] = pixel_val;
  assign array_175531[1] = pixel_val__1;
  assign array_175531[2] = pixel_val__2;
  assign array_175531[3] = pixel_val__3;
  assign out = {array_175531[3], array_175531[2], array_175531[1], array_175531[0]};
endmodule
