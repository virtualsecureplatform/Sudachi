module __riscv_simple__run_instruction(
  input wire [31:0] pc,
  input wire [31:0] ins,
  input wire [1023:0] regs,
  input wire [127:0] dmem,
  output wire [1183:0] out
);
  wire [31:0] regs_unflattened[32];
  assign regs_unflattened[0] = regs[31:0];
  assign regs_unflattened[1] = regs[63:32];
  assign regs_unflattened[2] = regs[95:64];
  assign regs_unflattened[3] = regs[127:96];
  assign regs_unflattened[4] = regs[159:128];
  assign regs_unflattened[5] = regs[191:160];
  assign regs_unflattened[6] = regs[223:192];
  assign regs_unflattened[7] = regs[255:224];
  assign regs_unflattened[8] = regs[287:256];
  assign regs_unflattened[9] = regs[319:288];
  assign regs_unflattened[10] = regs[351:320];
  assign regs_unflattened[11] = regs[383:352];
  assign regs_unflattened[12] = regs[415:384];
  assign regs_unflattened[13] = regs[447:416];
  assign regs_unflattened[14] = regs[479:448];
  assign regs_unflattened[15] = regs[511:480];
  assign regs_unflattened[16] = regs[543:512];
  assign regs_unflattened[17] = regs[575:544];
  assign regs_unflattened[18] = regs[607:576];
  assign regs_unflattened[19] = regs[639:608];
  assign regs_unflattened[20] = regs[671:640];
  assign regs_unflattened[21] = regs[703:672];
  assign regs_unflattened[22] = regs[735:704];
  assign regs_unflattened[23] = regs[767:736];
  assign regs_unflattened[24] = regs[799:768];
  assign regs_unflattened[25] = regs[831:800];
  assign regs_unflattened[26] = regs[863:832];
  assign regs_unflattened[27] = regs[895:864];
  assign regs_unflattened[28] = regs[927:896];
  assign regs_unflattened[29] = regs[959:928];
  assign regs_unflattened[30] = regs[991:960];
  assign regs_unflattened[31] = regs[1023:992];
  wire [7:0] dmem_unflattened[16];
  assign dmem_unflattened[0] = dmem[7:0];
  assign dmem_unflattened[1] = dmem[15:8];
  assign dmem_unflattened[2] = dmem[23:16];
  assign dmem_unflattened[3] = dmem[31:24];
  assign dmem_unflattened[4] = dmem[39:32];
  assign dmem_unflattened[5] = dmem[47:40];
  assign dmem_unflattened[6] = dmem[55:48];
  assign dmem_unflattened[7] = dmem[63:56];
  assign dmem_unflattened[8] = dmem[71:64];
  assign dmem_unflattened[9] = dmem[79:72];
  assign dmem_unflattened[10] = dmem[87:80];
  assign dmem_unflattened[11] = dmem[95:88];
  assign dmem_unflattened[12] = dmem[103:96];
  assign dmem_unflattened[13] = dmem[111:104];
  assign dmem_unflattened[14] = dmem[119:112];
  assign dmem_unflattened[15] = dmem[127:120];
  wire [4:0] rs1__5;
  wire [11:0] imm_11_0;
  wire [2:0] funct3__5;
  wire [2:0] ANDI;
  wire [2:0] ORI;
  wire [2:0] SRLI;
  wire [2:0] XORI;
  wire [2:0] SLLI;
  wire [2:0] ADDI;
  wire [31:0] array_index_3005;
  wire [31:0] concat_3006;
  wire eq_3007;
  wire eq_3008;
  wire eq_3009;
  wire eq_3010;
  wire eq_3011;
  wire eq_3012;
  wire [6:0] opcode__3;
  wire [6:0] I_LD__1;
  wire [2:0] LW;
  wire [31:0] addr;
  wire [6:0] I_ARITH__1;
  wire [6:0] I_JALR__1;
  wire [6:0] concat_3019;
  wire eq_3020;
  wire eq_3021;
  wire [6:0] R_CLASS;
  wire [6:0] S_CLASS;
  wire eq_3026;
  wire eq_3027;
  wire [6:0] B_CLASS;
  wire [6:0] U_CLASS;
  wire [6:0] UJ_CLASS;
  wire [7:0] one_hot_3031;
  wire [30:0] add_3034;
  wire imm_12;
  wire imm_11;
  wire [5:0] imm_10_5;
  wire [3:0] imm_4_1;
  wire [2:0] ADDI__1;
  wire eq_3041;
  wire eq_3042;
  wire or_3043;
  wire eq_3044;
  wire eq_3045;
  wire eq_3046;
  wire [6:0] funct7__1;
  wire [6:0] SRA_FUNCT7;
  wire [6:0] SRA_FUNCT7__1;
  wire [4:0] and_3053;
  wire [31:0] concat_3054;
  wire [4:0] rs2__1;
  wire [11:0] concat_3059;
  wire [6:0] and_3065;
  wire [7:0] array_index_3066;
  wire [31:0] add_3067;
  wire [7:0] array_index_3070;
  wire [31:0] add_3071;
  wire [29:0] add_3073;
  wire [2:0] LW__1;
  wire [4:0] rd__3;
  wire [31:0] array_index_3077;
  wire [7:0] imm_19_12;
  wire imm_11__1;
  wire [9:0] imm_10_1;
  wire [1:0] concat_3086;
  wire and_3088;
  wire [31:0] shll_3091;
  wire [31:0] xor_3092;
  wire [31:0] shrl_3093;
  wire [31:0] shra_3094;
  wire [31:0] or_3095;
  wire [31:0] sign_ext_3096;
  wire [7:0] array_index_3098;
  wire or_3100;
  wire [31:0] concat_3112;
  wire [30:0] add_3116;
  wire [19:0] concat_3118;
  wire or_3119;
  wire or_3120;
  wire [9:0] concat_3123;
  wire [9:0] concat_3134;
  wire [11:0] concat_3145;
  wire [31:0] add_3161;
  wire [31:0] add_3162;
  wire [30:0] add_3163;
  wire [31:0] new_rd;
  wire [31:0] pc_imm__2;
  wire or_3177;
  wire [7:0] concat_3178;
  wire [31:0] sub_3183;
  wire [31:0] add_3184;
  wire [19:0] imm_31_12;
  wire [6:0] S_CLASS__1;
  wire [3:0] and_3193;
  wire [7:0] dmem__3[16];
  wire [31:0] add_3196;
  wire [5:0] and_3199;
  wire [31:0] add_3200;
  wire [31:0] sel_3201;
  wire [31:0] sel_3202;
  wire [31:0] sel_3203;
  wire [31:0] sel_3204;
  wire [31:0] sel_3205;
  wire [31:0] sel_3206;
  wire [30:0] add_3207;
  wire [31:0] new_value;
  wire [31:0] new_value__1;
  wire [7:0] dmem__4[16];
  wire [31:0] add_3217;
  wire [31:0] add_3218;
  wire [9:0] concat_3222;
  wire [8:0] concat_3231;
  wire [6:0] concat_3241;
  wire [4:0] concat_3248;
  wire [31:0] array_update_3249[32];
  wire [31:0] array_update_3250[32];
  wire [31:0] array_update_3251[32];
  wire [31:0] array_update_3252[32];
  wire [7:0] dmem__5[16];
  wire [31:0] add_3257;
  wire [7:0] dmem__6[16];
  wire [31:0] regs__2[32];
  wire [3:0] concat_3268;
  wire [7:0] array_update_3269[16];
  wire [7:0] array_update_3270[16];
  wire [7:0] array_update_3271[16];
  wire [31:0] pc__3;
  wire [31:0] array_update_3277[32];
  wire [7:0] dmem__2[16];
  assign rs1__5 = ins[19:15];
  assign imm_11_0 = ins[31:20];
  assign funct3__5 = ins[14:12];
  assign ANDI = 3'h7;
  assign ORI = 3'h6;
  assign SRLI = 3'h5;
  assign XORI = 3'h4;
  assign SLLI = 3'h1;
  assign ADDI = 3'h0;
  assign array_index_3005 = regs_unflattened[rs1__5];
  assign concat_3006 = {20'h0_0000, imm_11_0};
  assign eq_3007 = funct3__5 == ANDI;
  assign eq_3008 = funct3__5 == ORI;
  assign eq_3009 = funct3__5 == SRLI;
  assign eq_3010 = funct3__5 == XORI;
  assign eq_3011 = funct3__5 == SLLI;
  assign eq_3012 = funct3__5 == ADDI;
  assign opcode__3 = ins[6:0];
  assign I_LD__1 = 7'h03;
  assign LW = 3'h2;
  assign addr = array_index_3005 + concat_3006;
  assign I_ARITH__1 = 7'h13;
  assign I_JALR__1 = 7'h67;
  assign concat_3019 = {eq_3007, eq_3008, eq_3009, eq_3009, eq_3010, eq_3011, eq_3012};
  assign eq_3020 = opcode__3 == I_LD__1;
  assign eq_3021 = funct3__5 == LW;
  assign R_CLASS = 7'h33;
  assign S_CLASS = 7'h23;
  assign eq_3026 = opcode__3 == I_ARITH__1;
  assign eq_3027 = opcode__3 == I_JALR__1;
  assign B_CLASS = 7'h63;
  assign U_CLASS = 7'h37;
  assign UJ_CLASS = 7'h6f;
  assign one_hot_3031 = {concat_3019[6:0] == 7'h00, concat_3019[6] && concat_3019[5:0] == 6'h00, concat_3019[5] && concat_3019[4:0] == 5'h00, concat_3019[4] && concat_3019[3:0] == 4'h0, concat_3019[3] && concat_3019[2:0] == 3'h0, concat_3019[2] && concat_3019[1:0] == 2'h0, concat_3019[1] && !concat_3019[0], concat_3019[0]};
  assign add_3034 = addr[31:1] + 31'h0000_0001;
  assign imm_12 = ins[31];
  assign imm_11 = ins[7];
  assign imm_10_5 = ins[30:25];
  assign imm_4_1 = ins[11:8];
  assign ADDI__1 = 3'h0;
  assign eq_3041 = opcode__3 == R_CLASS;
  assign eq_3042 = opcode__3 == S_CLASS;
  assign or_3043 = eq_3026 | eq_3027 | eq_3020;
  assign eq_3044 = opcode__3 == B_CLASS;
  assign eq_3045 = opcode__3 == U_CLASS;
  assign eq_3046 = opcode__3 == UJ_CLASS;
  assign funct7__1 = ins[31:25];
  assign SRA_FUNCT7 = 7'h20;
  assign SRA_FUNCT7__1 = 7'h20;
  assign and_3053 = {5{eq_3020}} & {eq_3009, eq_3010, eq_3021, eq_3011, eq_3012};
  assign concat_3054 = {add_3034, addr[0]};
  assign rs2__1 = ins[24:20];
  assign concat_3059 = {imm_12, imm_11, imm_10_5, imm_4_1};
  assign and_3065 = {7{eq_3026}} & one_hot_3031[6:0];
  assign array_index_3066 = dmem_unflattened[addr > 32'h0000_000f ? 4'hf : addr[3:0]];
  assign add_3067 = addr + 32'h0000_0001;
  assign array_index_3070 = dmem_unflattened[concat_3054 > 32'h0000_000f ? 4'hf : concat_3054[3:0]];
  assign add_3071 = addr + 32'h0000_0003;
  assign add_3073 = pc[31:2] + 30'h0000_0001;
  assign LW__1 = 3'h2;
  assign rd__3 = ins[11:7];
  assign array_index_3077 = regs_unflattened[rs2__1];
  assign imm_19_12 = ins[19:12];
  assign imm_11__1 = ins[20];
  assign imm_10_1 = ins[30:21];
  assign concat_3086 = {funct7__1 != SRA_FUNCT7, funct7__1 == SRA_FUNCT7__1};
  assign and_3088 = eq_3027 & eq_3012;
  assign shll_3091 = imm_11_0 >= 12'h020 ? 32'h0000_0000 : array_index_3005 << imm_11_0;
  assign xor_3092 = array_index_3005 ^ concat_3006;
  assign shrl_3093 = imm_11_0 >= 12'h020 ? 32'h0000_0000 : array_index_3005 >> imm_11_0;
  assign shra_3094 = imm_11_0 >= 12'h020 ? {32{array_index_3005[31]}} : $unsigned($signed(array_index_3005) >>> imm_11_0);
  assign or_3095 = array_index_3005 | concat_3006;
  assign sign_ext_3096 = {{24{array_index_3066[7]}}, array_index_3066};
  assign array_index_3098 = dmem_unflattened[add_3067 > 32'h0000_000f ? 4'hf : add_3067[3:0]];
  assign or_3100 = and_3053[1] | and_3053[4];
  assign concat_3112 = {20'h0_0000, funct7__1, rd__3};
  assign add_3116 = pc[31:1] + {{19{concat_3059[11]}}, concat_3059};
  assign concat_3118 = {imm_12, imm_19_12, imm_11__1, imm_10_1};
  assign or_3119 = eq_3041 | eq_3042 | eq_3045 | eq_3026 | eq_3020;
  assign or_3120 = or_3043 & ~(eq_3026 | eq_3020) & eq_3027 & funct3__5 != ADDI__1 | ~(eq_3041 | eq_3042 | or_3043 | eq_3044 | eq_3045 | eq_3046);
  assign concat_3123 = {and_3088, and_3053[2:0], and_3065[5:0]};
  assign concat_3134 = {and_3088, and_3053[2], or_3100, and_3053[0], and_3065[5:0]};
  assign concat_3145 = {and_3088, and_3053[3:2], or_3100, and_3053[0], and_3065};
  assign add_3161 = array_index_3077 + concat_3112;
  assign add_3162 = array_index_3077 + 32'h0000_0001;
  assign add_3163 = array_index_3077[31:1] + 31'h0000_0001;
  assign new_rd = {add_3073, pc[1:0]};
  assign pc_imm__2 = {add_3116, pc[0]};
  assign or_3177 = or_3119 | or_3120;
  assign concat_3178 = {{2{eq_3009}} & concat_3086, {2{eq_3012}} & concat_3086, eq_3011, eq_3008, eq_3007, eq_3010};
  assign sub_3183 = array_index_3005 - array_index_3077;
  assign add_3184 = array_index_3005 + array_index_3077;
  assign imm_31_12 = ins[31:12];
  assign S_CLASS__1 = 7'h23;
  assign and_3193 = {4{eq_3042}} & {funct3__5 > LW__1, eq_3012, eq_3011, eq_3021};
  assign dmem__3[0] = add_3161 == 32'h0000_0000 ? array_index_3005[31:24] : dmem_unflattened[0];
  assign dmem__3[1] = add_3161 == 32'h0000_0001 ? array_index_3005[31:24] : dmem_unflattened[1];
  assign dmem__3[2] = add_3161 == 32'h0000_0002 ? array_index_3005[31:24] : dmem_unflattened[2];
  assign dmem__3[3] = add_3161 == 32'h0000_0003 ? array_index_3005[31:24] : dmem_unflattened[3];
  assign dmem__3[4] = add_3161 == 32'h0000_0004 ? array_index_3005[31:24] : dmem_unflattened[4];
  assign dmem__3[5] = add_3161 == 32'h0000_0005 ? array_index_3005[31:24] : dmem_unflattened[5];
  assign dmem__3[6] = add_3161 == 32'h0000_0006 ? array_index_3005[31:24] : dmem_unflattened[6];
  assign dmem__3[7] = add_3161 == 32'h0000_0007 ? array_index_3005[31:24] : dmem_unflattened[7];
  assign dmem__3[8] = add_3161 == 32'h0000_0008 ? array_index_3005[31:24] : dmem_unflattened[8];
  assign dmem__3[9] = add_3161 == 32'h0000_0009 ? array_index_3005[31:24] : dmem_unflattened[9];
  assign dmem__3[10] = add_3161 == 32'h0000_000a ? array_index_3005[31:24] : dmem_unflattened[10];
  assign dmem__3[11] = add_3161 == 32'h0000_000b ? array_index_3005[31:24] : dmem_unflattened[11];
  assign dmem__3[12] = add_3161 == 32'h0000_000c ? array_index_3005[31:24] : dmem_unflattened[12];
  assign dmem__3[13] = add_3161 == 32'h0000_000d ? array_index_3005[31:24] : dmem_unflattened[13];
  assign dmem__3[14] = add_3161 == 32'h0000_000e ? array_index_3005[31:24] : dmem_unflattened[14];
  assign dmem__3[15] = add_3161 == 32'h0000_000f ? array_index_3005[31:24] : dmem_unflattened[15];
  assign add_3196 = add_3162 + concat_3112;
  assign and_3199 = {6{eq_3044}} & {eq_3007, eq_3008, eq_3009, eq_3010, eq_3011, eq_3012};
  assign add_3200 = array_index_3005 + {{20{imm_11_0[11]}}, imm_11_0};
  assign sel_3201 = array_index_3005 == array_index_3077 ? pc_imm__2 : new_rd;
  assign sel_3202 = array_index_3005 != array_index_3077 ? pc_imm__2 : new_rd;
  assign sel_3203 = $signed(array_index_3005) < $signed(array_index_3077) ? pc_imm__2 : new_rd;
  assign sel_3204 = $signed(array_index_3005) >= $signed(array_index_3077) ? pc_imm__2 : new_rd;
  assign sel_3205 = array_index_3005 < array_index_3077 ? pc_imm__2 : new_rd;
  assign sel_3206 = array_index_3005 >= array_index_3077 ? pc_imm__2 : new_rd;
  assign add_3207 = pc[31:1] + {{11{concat_3118[19]}}, concat_3118};
  assign new_value = (array_index_3005 ^ array_index_3077) & {32{concat_3178[0]}} | array_index_3005 & array_index_3077 & {32{concat_3178[1]}} | (array_index_3005 | array_index_3077) & {32{concat_3178[2]}} | (array_index_3077 >= 32'h0000_0020 ? 32'h0000_0000 : array_index_3005 << array_index_3077) & {32{concat_3178[3]}} | sub_3183 & {32{concat_3178[4]}} | add_3184 & {32{concat_3178[5]}} | (array_index_3077 >= 32'h0000_0020 ? {32{array_index_3005[31]}} : $unsigned($signed(array_index_3005) >>> array_index_3077)) & {32{concat_3178[6]}} | (array_index_3077 >= 32'h0000_0020 ? 32'h0000_0000 : array_index_3005 >> array_index_3077) & {32{concat_3178[7]}};
  assign new_value__1 = {addr[31:16] & {16{concat_3123[0]}} | shll_3091[31:16] & {16{concat_3123[1]}} | xor_3092[31:16] & {16{concat_3123[2]}} | shrl_3093[31:16] & {16{concat_3123[3]}} | shra_3094[31:16] & {16{concat_3123[4]}} | or_3095[31:16] & {16{concat_3123[5]}} | sign_ext_3096[31:16] & {16{concat_3123[6]}} | {16{array_index_3066[7]}} & {16{concat_3123[7]}} | {array_index_3066, array_index_3098} & {16{concat_3123[8]}} | add_3073[29:14] & {16{concat_3123[9]}}, addr[15:12] & {4{concat_3134[0]}} | shll_3091[15:12] & {4{concat_3134[1]}} | xor_3092[15:12] & {4{concat_3134[2]}} | shrl_3093[15:12] & {4{concat_3134[3]}} | shra_3094[15:12] & {4{concat_3134[4]}} | or_3095[15:12] & {4{concat_3134[5]}} | sign_ext_3096[15:12] & {4{concat_3134[6]}} | array_index_3066[7:4] & {4{concat_3134[7]}} | array_index_3070[7:4] & {4{concat_3134[8]}} | add_3073[13:10] & {4{concat_3134[9]}}, addr[11:0] & {12{concat_3145[0]}} | shll_3091[11:0] & {12{concat_3145[1]}} | xor_3092[11:0] & {12{concat_3145[2]}} | shrl_3093[11:0] & {12{concat_3145[3]}} | shra_3094[11:0] & {12{concat_3145[4]}} | or_3095[11:0] & {12{concat_3145[5]}} | array_index_3005[11:0] & imm_11_0 & {12{concat_3145[6]}} | sign_ext_3096[11:0] & {12{concat_3145[7]}} | {array_index_3066[3:0], array_index_3098} & {12{concat_3145[8]}} | {array_index_3070[3:0], dmem_unflattened[add_3071 > 32'h0000_000f ? 4'hf : add_3071[3:0]]} & {12{concat_3145[9]}} | {4'h0, dmem_unflattened[regs_unflattened[addr > 32'h0000_001f ? 5'h1f : addr[4:0]] > 32'h0000_000f ? 4'hf : regs_unflattened[addr > 32'h0000_001f ? 5'h1f : addr[4:0]][3:0]]} & {12{concat_3145[10]}} | {add_3073[9:0], pc[1:0]} & {12{concat_3145[11]}}};
  assign dmem__4[0] = add_3196 == 32'h0000_0000 ? array_index_3005[23:16] : dmem__3[0];
  assign dmem__4[1] = add_3196 == 32'h0000_0001 ? array_index_3005[23:16] : dmem__3[1];
  assign dmem__4[2] = add_3196 == 32'h0000_0002 ? array_index_3005[23:16] : dmem__3[2];
  assign dmem__4[3] = add_3196 == 32'h0000_0003 ? array_index_3005[23:16] : dmem__3[3];
  assign dmem__4[4] = add_3196 == 32'h0000_0004 ? array_index_3005[23:16] : dmem__3[4];
  assign dmem__4[5] = add_3196 == 32'h0000_0005 ? array_index_3005[23:16] : dmem__3[5];
  assign dmem__4[6] = add_3196 == 32'h0000_0006 ? array_index_3005[23:16] : dmem__3[6];
  assign dmem__4[7] = add_3196 == 32'h0000_0007 ? array_index_3005[23:16] : dmem__3[7];
  assign dmem__4[8] = add_3196 == 32'h0000_0008 ? array_index_3005[23:16] : dmem__3[8];
  assign dmem__4[9] = add_3196 == 32'h0000_0009 ? array_index_3005[23:16] : dmem__3[9];
  assign dmem__4[10] = add_3196 == 32'h0000_000a ? array_index_3005[23:16] : dmem__3[10];
  assign dmem__4[11] = add_3196 == 32'h0000_000b ? array_index_3005[23:16] : dmem__3[11];
  assign dmem__4[12] = add_3196 == 32'h0000_000c ? array_index_3005[23:16] : dmem__3[12];
  assign dmem__4[13] = add_3196 == 32'h0000_000d ? array_index_3005[23:16] : dmem__3[13];
  assign dmem__4[14] = add_3196 == 32'h0000_000e ? array_index_3005[23:16] : dmem__3[14];
  assign dmem__4[15] = add_3196 == 32'h0000_000f ? array_index_3005[23:16] : dmem__3[15];
  assign add_3217 = {add_3163, array_index_3077[0]} + concat_3112;
  assign add_3218 = array_index_3077 + 32'h0000_0003;
  assign concat_3222 = {eq_3046, and_3199, or_3120, and_3088, or_3119};
  assign concat_3231 = {eq_3046, and_3199, and_3088, or_3177};
  assign concat_3241 = {and_3199, or_3177 | eq_3046};
  assign concat_3248 = {eq_3046, eq_3045, or_3043, eq_3042 | eq_3044 | ~(eq_3041 | eq_3042 | or_3043 | eq_3044 | eq_3045 | eq_3046), eq_3041};
  assign array_update_3249[0] = rd__3 == 5'h00 ? new_value : regs_unflattened[0];
  assign array_update_3249[1] = rd__3 == 5'h01 ? new_value : regs_unflattened[1];
  assign array_update_3249[2] = rd__3 == 5'h02 ? new_value : regs_unflattened[2];
  assign array_update_3249[3] = rd__3 == 5'h03 ? new_value : regs_unflattened[3];
  assign array_update_3249[4] = rd__3 == 5'h04 ? new_value : regs_unflattened[4];
  assign array_update_3249[5] = rd__3 == 5'h05 ? new_value : regs_unflattened[5];
  assign array_update_3249[6] = rd__3 == 5'h06 ? new_value : regs_unflattened[6];
  assign array_update_3249[7] = rd__3 == 5'h07 ? new_value : regs_unflattened[7];
  assign array_update_3249[8] = rd__3 == 5'h08 ? new_value : regs_unflattened[8];
  assign array_update_3249[9] = rd__3 == 5'h09 ? new_value : regs_unflattened[9];
  assign array_update_3249[10] = rd__3 == 5'h0a ? new_value : regs_unflattened[10];
  assign array_update_3249[11] = rd__3 == 5'h0b ? new_value : regs_unflattened[11];
  assign array_update_3249[12] = rd__3 == 5'h0c ? new_value : regs_unflattened[12];
  assign array_update_3249[13] = rd__3 == 5'h0d ? new_value : regs_unflattened[13];
  assign array_update_3249[14] = rd__3 == 5'h0e ? new_value : regs_unflattened[14];
  assign array_update_3249[15] = rd__3 == 5'h0f ? new_value : regs_unflattened[15];
  assign array_update_3249[16] = rd__3 == 5'h10 ? new_value : regs_unflattened[16];
  assign array_update_3249[17] = rd__3 == 5'h11 ? new_value : regs_unflattened[17];
  assign array_update_3249[18] = rd__3 == 5'h12 ? new_value : regs_unflattened[18];
  assign array_update_3249[19] = rd__3 == 5'h13 ? new_value : regs_unflattened[19];
  assign array_update_3249[20] = rd__3 == 5'h14 ? new_value : regs_unflattened[20];
  assign array_update_3249[21] = rd__3 == 5'h15 ? new_value : regs_unflattened[21];
  assign array_update_3249[22] = rd__3 == 5'h16 ? new_value : regs_unflattened[22];
  assign array_update_3249[23] = rd__3 == 5'h17 ? new_value : regs_unflattened[23];
  assign array_update_3249[24] = rd__3 == 5'h18 ? new_value : regs_unflattened[24];
  assign array_update_3249[25] = rd__3 == 5'h19 ? new_value : regs_unflattened[25];
  assign array_update_3249[26] = rd__3 == 5'h1a ? new_value : regs_unflattened[26];
  assign array_update_3249[27] = rd__3 == 5'h1b ? new_value : regs_unflattened[27];
  assign array_update_3249[28] = rd__3 == 5'h1c ? new_value : regs_unflattened[28];
  assign array_update_3249[29] = rd__3 == 5'h1d ? new_value : regs_unflattened[29];
  assign array_update_3249[30] = rd__3 == 5'h1e ? new_value : regs_unflattened[30];
  assign array_update_3249[31] = rd__3 == 5'h1f ? new_value : regs_unflattened[31];
  assign array_update_3250[0] = rd__3 == 5'h00 ? new_value__1 : regs_unflattened[0];
  assign array_update_3250[1] = rd__3 == 5'h01 ? new_value__1 : regs_unflattened[1];
  assign array_update_3250[2] = rd__3 == 5'h02 ? new_value__1 : regs_unflattened[2];
  assign array_update_3250[3] = rd__3 == 5'h03 ? new_value__1 : regs_unflattened[3];
  assign array_update_3250[4] = rd__3 == 5'h04 ? new_value__1 : regs_unflattened[4];
  assign array_update_3250[5] = rd__3 == 5'h05 ? new_value__1 : regs_unflattened[5];
  assign array_update_3250[6] = rd__3 == 5'h06 ? new_value__1 : regs_unflattened[6];
  assign array_update_3250[7] = rd__3 == 5'h07 ? new_value__1 : regs_unflattened[7];
  assign array_update_3250[8] = rd__3 == 5'h08 ? new_value__1 : regs_unflattened[8];
  assign array_update_3250[9] = rd__3 == 5'h09 ? new_value__1 : regs_unflattened[9];
  assign array_update_3250[10] = rd__3 == 5'h0a ? new_value__1 : regs_unflattened[10];
  assign array_update_3250[11] = rd__3 == 5'h0b ? new_value__1 : regs_unflattened[11];
  assign array_update_3250[12] = rd__3 == 5'h0c ? new_value__1 : regs_unflattened[12];
  assign array_update_3250[13] = rd__3 == 5'h0d ? new_value__1 : regs_unflattened[13];
  assign array_update_3250[14] = rd__3 == 5'h0e ? new_value__1 : regs_unflattened[14];
  assign array_update_3250[15] = rd__3 == 5'h0f ? new_value__1 : regs_unflattened[15];
  assign array_update_3250[16] = rd__3 == 5'h10 ? new_value__1 : regs_unflattened[16];
  assign array_update_3250[17] = rd__3 == 5'h11 ? new_value__1 : regs_unflattened[17];
  assign array_update_3250[18] = rd__3 == 5'h12 ? new_value__1 : regs_unflattened[18];
  assign array_update_3250[19] = rd__3 == 5'h13 ? new_value__1 : regs_unflattened[19];
  assign array_update_3250[20] = rd__3 == 5'h14 ? new_value__1 : regs_unflattened[20];
  assign array_update_3250[21] = rd__3 == 5'h15 ? new_value__1 : regs_unflattened[21];
  assign array_update_3250[22] = rd__3 == 5'h16 ? new_value__1 : regs_unflattened[22];
  assign array_update_3250[23] = rd__3 == 5'h17 ? new_value__1 : regs_unflattened[23];
  assign array_update_3250[24] = rd__3 == 5'h18 ? new_value__1 : regs_unflattened[24];
  assign array_update_3250[25] = rd__3 == 5'h19 ? new_value__1 : regs_unflattened[25];
  assign array_update_3250[26] = rd__3 == 5'h1a ? new_value__1 : regs_unflattened[26];
  assign array_update_3250[27] = rd__3 == 5'h1b ? new_value__1 : regs_unflattened[27];
  assign array_update_3250[28] = rd__3 == 5'h1c ? new_value__1 : regs_unflattened[28];
  assign array_update_3250[29] = rd__3 == 5'h1d ? new_value__1 : regs_unflattened[29];
  assign array_update_3250[30] = rd__3 == 5'h1e ? new_value__1 : regs_unflattened[30];
  assign array_update_3250[31] = rd__3 == 5'h1f ? new_value__1 : regs_unflattened[31];
  assign array_update_3251[0] = rd__3 == 5'h00 ? {imm_31_12, 12'h000} : regs_unflattened[0];
  assign array_update_3251[1] = rd__3 == 5'h01 ? {imm_31_12, 12'h000} : regs_unflattened[1];
  assign array_update_3251[2] = rd__3 == 5'h02 ? {imm_31_12, 12'h000} : regs_unflattened[2];
  assign array_update_3251[3] = rd__3 == 5'h03 ? {imm_31_12, 12'h000} : regs_unflattened[3];
  assign array_update_3251[4] = rd__3 == 5'h04 ? {imm_31_12, 12'h000} : regs_unflattened[4];
  assign array_update_3251[5] = rd__3 == 5'h05 ? {imm_31_12, 12'h000} : regs_unflattened[5];
  assign array_update_3251[6] = rd__3 == 5'h06 ? {imm_31_12, 12'h000} : regs_unflattened[6];
  assign array_update_3251[7] = rd__3 == 5'h07 ? {imm_31_12, 12'h000} : regs_unflattened[7];
  assign array_update_3251[8] = rd__3 == 5'h08 ? {imm_31_12, 12'h000} : regs_unflattened[8];
  assign array_update_3251[9] = rd__3 == 5'h09 ? {imm_31_12, 12'h000} : regs_unflattened[9];
  assign array_update_3251[10] = rd__3 == 5'h0a ? {imm_31_12, 12'h000} : regs_unflattened[10];
  assign array_update_3251[11] = rd__3 == 5'h0b ? {imm_31_12, 12'h000} : regs_unflattened[11];
  assign array_update_3251[12] = rd__3 == 5'h0c ? {imm_31_12, 12'h000} : regs_unflattened[12];
  assign array_update_3251[13] = rd__3 == 5'h0d ? {imm_31_12, 12'h000} : regs_unflattened[13];
  assign array_update_3251[14] = rd__3 == 5'h0e ? {imm_31_12, 12'h000} : regs_unflattened[14];
  assign array_update_3251[15] = rd__3 == 5'h0f ? {imm_31_12, 12'h000} : regs_unflattened[15];
  assign array_update_3251[16] = rd__3 == 5'h10 ? {imm_31_12, 12'h000} : regs_unflattened[16];
  assign array_update_3251[17] = rd__3 == 5'h11 ? {imm_31_12, 12'h000} : regs_unflattened[17];
  assign array_update_3251[18] = rd__3 == 5'h12 ? {imm_31_12, 12'h000} : regs_unflattened[18];
  assign array_update_3251[19] = rd__3 == 5'h13 ? {imm_31_12, 12'h000} : regs_unflattened[19];
  assign array_update_3251[20] = rd__3 == 5'h14 ? {imm_31_12, 12'h000} : regs_unflattened[20];
  assign array_update_3251[21] = rd__3 == 5'h15 ? {imm_31_12, 12'h000} : regs_unflattened[21];
  assign array_update_3251[22] = rd__3 == 5'h16 ? {imm_31_12, 12'h000} : regs_unflattened[22];
  assign array_update_3251[23] = rd__3 == 5'h17 ? {imm_31_12, 12'h000} : regs_unflattened[23];
  assign array_update_3251[24] = rd__3 == 5'h18 ? {imm_31_12, 12'h000} : regs_unflattened[24];
  assign array_update_3251[25] = rd__3 == 5'h19 ? {imm_31_12, 12'h000} : regs_unflattened[25];
  assign array_update_3251[26] = rd__3 == 5'h1a ? {imm_31_12, 12'h000} : regs_unflattened[26];
  assign array_update_3251[27] = rd__3 == 5'h1b ? {imm_31_12, 12'h000} : regs_unflattened[27];
  assign array_update_3251[28] = rd__3 == 5'h1c ? {imm_31_12, 12'h000} : regs_unflattened[28];
  assign array_update_3251[29] = rd__3 == 5'h1d ? {imm_31_12, 12'h000} : regs_unflattened[29];
  assign array_update_3251[30] = rd__3 == 5'h1e ? {imm_31_12, 12'h000} : regs_unflattened[30];
  assign array_update_3251[31] = rd__3 == 5'h1f ? {imm_31_12, 12'h000} : regs_unflattened[31];
  assign array_update_3252[0] = rd__3 == 5'h00 ? new_rd : regs_unflattened[0];
  assign array_update_3252[1] = rd__3 == 5'h01 ? new_rd : regs_unflattened[1];
  assign array_update_3252[2] = rd__3 == 5'h02 ? new_rd : regs_unflattened[2];
  assign array_update_3252[3] = rd__3 == 5'h03 ? new_rd : regs_unflattened[3];
  assign array_update_3252[4] = rd__3 == 5'h04 ? new_rd : regs_unflattened[4];
  assign array_update_3252[5] = rd__3 == 5'h05 ? new_rd : regs_unflattened[5];
  assign array_update_3252[6] = rd__3 == 5'h06 ? new_rd : regs_unflattened[6];
  assign array_update_3252[7] = rd__3 == 5'h07 ? new_rd : regs_unflattened[7];
  assign array_update_3252[8] = rd__3 == 5'h08 ? new_rd : regs_unflattened[8];
  assign array_update_3252[9] = rd__3 == 5'h09 ? new_rd : regs_unflattened[9];
  assign array_update_3252[10] = rd__3 == 5'h0a ? new_rd : regs_unflattened[10];
  assign array_update_3252[11] = rd__3 == 5'h0b ? new_rd : regs_unflattened[11];
  assign array_update_3252[12] = rd__3 == 5'h0c ? new_rd : regs_unflattened[12];
  assign array_update_3252[13] = rd__3 == 5'h0d ? new_rd : regs_unflattened[13];
  assign array_update_3252[14] = rd__3 == 5'h0e ? new_rd : regs_unflattened[14];
  assign array_update_3252[15] = rd__3 == 5'h0f ? new_rd : regs_unflattened[15];
  assign array_update_3252[16] = rd__3 == 5'h10 ? new_rd : regs_unflattened[16];
  assign array_update_3252[17] = rd__3 == 5'h11 ? new_rd : regs_unflattened[17];
  assign array_update_3252[18] = rd__3 == 5'h12 ? new_rd : regs_unflattened[18];
  assign array_update_3252[19] = rd__3 == 5'h13 ? new_rd : regs_unflattened[19];
  assign array_update_3252[20] = rd__3 == 5'h14 ? new_rd : regs_unflattened[20];
  assign array_update_3252[21] = rd__3 == 5'h15 ? new_rd : regs_unflattened[21];
  assign array_update_3252[22] = rd__3 == 5'h16 ? new_rd : regs_unflattened[22];
  assign array_update_3252[23] = rd__3 == 5'h17 ? new_rd : regs_unflattened[23];
  assign array_update_3252[24] = rd__3 == 5'h18 ? new_rd : regs_unflattened[24];
  assign array_update_3252[25] = rd__3 == 5'h19 ? new_rd : regs_unflattened[25];
  assign array_update_3252[26] = rd__3 == 5'h1a ? new_rd : regs_unflattened[26];
  assign array_update_3252[27] = rd__3 == 5'h1b ? new_rd : regs_unflattened[27];
  assign array_update_3252[28] = rd__3 == 5'h1c ? new_rd : regs_unflattened[28];
  assign array_update_3252[29] = rd__3 == 5'h1d ? new_rd : regs_unflattened[29];
  assign array_update_3252[30] = rd__3 == 5'h1e ? new_rd : regs_unflattened[30];
  assign array_update_3252[31] = rd__3 == 5'h1f ? new_rd : regs_unflattened[31];
  assign dmem__5[0] = add_3217 == 32'h0000_0000 ? array_index_3005[15:8] : dmem__4[0];
  assign dmem__5[1] = add_3217 == 32'h0000_0001 ? array_index_3005[15:8] : dmem__4[1];
  assign dmem__5[2] = add_3217 == 32'h0000_0002 ? array_index_3005[15:8] : dmem__4[2];
  assign dmem__5[3] = add_3217 == 32'h0000_0003 ? array_index_3005[15:8] : dmem__4[3];
  assign dmem__5[4] = add_3217 == 32'h0000_0004 ? array_index_3005[15:8] : dmem__4[4];
  assign dmem__5[5] = add_3217 == 32'h0000_0005 ? array_index_3005[15:8] : dmem__4[5];
  assign dmem__5[6] = add_3217 == 32'h0000_0006 ? array_index_3005[15:8] : dmem__4[6];
  assign dmem__5[7] = add_3217 == 32'h0000_0007 ? array_index_3005[15:8] : dmem__4[7];
  assign dmem__5[8] = add_3217 == 32'h0000_0008 ? array_index_3005[15:8] : dmem__4[8];
  assign dmem__5[9] = add_3217 == 32'h0000_0009 ? array_index_3005[15:8] : dmem__4[9];
  assign dmem__5[10] = add_3217 == 32'h0000_000a ? array_index_3005[15:8] : dmem__4[10];
  assign dmem__5[11] = add_3217 == 32'h0000_000b ? array_index_3005[15:8] : dmem__4[11];
  assign dmem__5[12] = add_3217 == 32'h0000_000c ? array_index_3005[15:8] : dmem__4[12];
  assign dmem__5[13] = add_3217 == 32'h0000_000d ? array_index_3005[15:8] : dmem__4[13];
  assign dmem__5[14] = add_3217 == 32'h0000_000e ? array_index_3005[15:8] : dmem__4[14];
  assign dmem__5[15] = add_3217 == 32'h0000_000f ? array_index_3005[15:8] : dmem__4[15];
  assign add_3257 = add_3218 + concat_3112;
  assign dmem__6[0] = add_3161 == 32'h0000_0000 ? array_index_3005[15:8] : dmem_unflattened[0];
  assign dmem__6[1] = add_3161 == 32'h0000_0001 ? array_index_3005[15:8] : dmem_unflattened[1];
  assign dmem__6[2] = add_3161 == 32'h0000_0002 ? array_index_3005[15:8] : dmem_unflattened[2];
  assign dmem__6[3] = add_3161 == 32'h0000_0003 ? array_index_3005[15:8] : dmem_unflattened[3];
  assign dmem__6[4] = add_3161 == 32'h0000_0004 ? array_index_3005[15:8] : dmem_unflattened[4];
  assign dmem__6[5] = add_3161 == 32'h0000_0005 ? array_index_3005[15:8] : dmem_unflattened[5];
  assign dmem__6[6] = add_3161 == 32'h0000_0006 ? array_index_3005[15:8] : dmem_unflattened[6];
  assign dmem__6[7] = add_3161 == 32'h0000_0007 ? array_index_3005[15:8] : dmem_unflattened[7];
  assign dmem__6[8] = add_3161 == 32'h0000_0008 ? array_index_3005[15:8] : dmem_unflattened[8];
  assign dmem__6[9] = add_3161 == 32'h0000_0009 ? array_index_3005[15:8] : dmem_unflattened[9];
  assign dmem__6[10] = add_3161 == 32'h0000_000a ? array_index_3005[15:8] : dmem_unflattened[10];
  assign dmem__6[11] = add_3161 == 32'h0000_000b ? array_index_3005[15:8] : dmem_unflattened[11];
  assign dmem__6[12] = add_3161 == 32'h0000_000c ? array_index_3005[15:8] : dmem_unflattened[12];
  assign dmem__6[13] = add_3161 == 32'h0000_000d ? array_index_3005[15:8] : dmem_unflattened[13];
  assign dmem__6[14] = add_3161 == 32'h0000_000e ? array_index_3005[15:8] : dmem_unflattened[14];
  assign dmem__6[15] = add_3161 == 32'h0000_000f ? array_index_3005[15:8] : dmem_unflattened[15];
  assign regs__2[0] = array_update_3249[0] & {32{concat_3248[0]}} | regs_unflattened[0] & {32{concat_3248[1]}} | array_update_3250[0] & {32{concat_3248[2]}} | array_update_3251[0] & {32{concat_3248[3]}} | array_update_3252[0] & {32{concat_3248[4]}};
  assign regs__2[1] = array_update_3249[1] & {32{concat_3248[0]}} | regs_unflattened[1] & {32{concat_3248[1]}} | array_update_3250[1] & {32{concat_3248[2]}} | array_update_3251[1] & {32{concat_3248[3]}} | array_update_3252[1] & {32{concat_3248[4]}};
  assign regs__2[2] = array_update_3249[2] & {32{concat_3248[0]}} | regs_unflattened[2] & {32{concat_3248[1]}} | array_update_3250[2] & {32{concat_3248[2]}} | array_update_3251[2] & {32{concat_3248[3]}} | array_update_3252[2] & {32{concat_3248[4]}};
  assign regs__2[3] = array_update_3249[3] & {32{concat_3248[0]}} | regs_unflattened[3] & {32{concat_3248[1]}} | array_update_3250[3] & {32{concat_3248[2]}} | array_update_3251[3] & {32{concat_3248[3]}} | array_update_3252[3] & {32{concat_3248[4]}};
  assign regs__2[4] = array_update_3249[4] & {32{concat_3248[0]}} | regs_unflattened[4] & {32{concat_3248[1]}} | array_update_3250[4] & {32{concat_3248[2]}} | array_update_3251[4] & {32{concat_3248[3]}} | array_update_3252[4] & {32{concat_3248[4]}};
  assign regs__2[5] = array_update_3249[5] & {32{concat_3248[0]}} | regs_unflattened[5] & {32{concat_3248[1]}} | array_update_3250[5] & {32{concat_3248[2]}} | array_update_3251[5] & {32{concat_3248[3]}} | array_update_3252[5] & {32{concat_3248[4]}};
  assign regs__2[6] = array_update_3249[6] & {32{concat_3248[0]}} | regs_unflattened[6] & {32{concat_3248[1]}} | array_update_3250[6] & {32{concat_3248[2]}} | array_update_3251[6] & {32{concat_3248[3]}} | array_update_3252[6] & {32{concat_3248[4]}};
  assign regs__2[7] = array_update_3249[7] & {32{concat_3248[0]}} | regs_unflattened[7] & {32{concat_3248[1]}} | array_update_3250[7] & {32{concat_3248[2]}} | array_update_3251[7] & {32{concat_3248[3]}} | array_update_3252[7] & {32{concat_3248[4]}};
  assign regs__2[8] = array_update_3249[8] & {32{concat_3248[0]}} | regs_unflattened[8] & {32{concat_3248[1]}} | array_update_3250[8] & {32{concat_3248[2]}} | array_update_3251[8] & {32{concat_3248[3]}} | array_update_3252[8] & {32{concat_3248[4]}};
  assign regs__2[9] = array_update_3249[9] & {32{concat_3248[0]}} | regs_unflattened[9] & {32{concat_3248[1]}} | array_update_3250[9] & {32{concat_3248[2]}} | array_update_3251[9] & {32{concat_3248[3]}} | array_update_3252[9] & {32{concat_3248[4]}};
  assign regs__2[10] = array_update_3249[10] & {32{concat_3248[0]}} | regs_unflattened[10] & {32{concat_3248[1]}} | array_update_3250[10] & {32{concat_3248[2]}} | array_update_3251[10] & {32{concat_3248[3]}} | array_update_3252[10] & {32{concat_3248[4]}};
  assign regs__2[11] = array_update_3249[11] & {32{concat_3248[0]}} | regs_unflattened[11] & {32{concat_3248[1]}} | array_update_3250[11] & {32{concat_3248[2]}} | array_update_3251[11] & {32{concat_3248[3]}} | array_update_3252[11] & {32{concat_3248[4]}};
  assign regs__2[12] = array_update_3249[12] & {32{concat_3248[0]}} | regs_unflattened[12] & {32{concat_3248[1]}} | array_update_3250[12] & {32{concat_3248[2]}} | array_update_3251[12] & {32{concat_3248[3]}} | array_update_3252[12] & {32{concat_3248[4]}};
  assign regs__2[13] = array_update_3249[13] & {32{concat_3248[0]}} | regs_unflattened[13] & {32{concat_3248[1]}} | array_update_3250[13] & {32{concat_3248[2]}} | array_update_3251[13] & {32{concat_3248[3]}} | array_update_3252[13] & {32{concat_3248[4]}};
  assign regs__2[14] = array_update_3249[14] & {32{concat_3248[0]}} | regs_unflattened[14] & {32{concat_3248[1]}} | array_update_3250[14] & {32{concat_3248[2]}} | array_update_3251[14] & {32{concat_3248[3]}} | array_update_3252[14] & {32{concat_3248[4]}};
  assign regs__2[15] = array_update_3249[15] & {32{concat_3248[0]}} | regs_unflattened[15] & {32{concat_3248[1]}} | array_update_3250[15] & {32{concat_3248[2]}} | array_update_3251[15] & {32{concat_3248[3]}} | array_update_3252[15] & {32{concat_3248[4]}};
  assign regs__2[16] = array_update_3249[16] & {32{concat_3248[0]}} | regs_unflattened[16] & {32{concat_3248[1]}} | array_update_3250[16] & {32{concat_3248[2]}} | array_update_3251[16] & {32{concat_3248[3]}} | array_update_3252[16] & {32{concat_3248[4]}};
  assign regs__2[17] = array_update_3249[17] & {32{concat_3248[0]}} | regs_unflattened[17] & {32{concat_3248[1]}} | array_update_3250[17] & {32{concat_3248[2]}} | array_update_3251[17] & {32{concat_3248[3]}} | array_update_3252[17] & {32{concat_3248[4]}};
  assign regs__2[18] = array_update_3249[18] & {32{concat_3248[0]}} | regs_unflattened[18] & {32{concat_3248[1]}} | array_update_3250[18] & {32{concat_3248[2]}} | array_update_3251[18] & {32{concat_3248[3]}} | array_update_3252[18] & {32{concat_3248[4]}};
  assign regs__2[19] = array_update_3249[19] & {32{concat_3248[0]}} | regs_unflattened[19] & {32{concat_3248[1]}} | array_update_3250[19] & {32{concat_3248[2]}} | array_update_3251[19] & {32{concat_3248[3]}} | array_update_3252[19] & {32{concat_3248[4]}};
  assign regs__2[20] = array_update_3249[20] & {32{concat_3248[0]}} | regs_unflattened[20] & {32{concat_3248[1]}} | array_update_3250[20] & {32{concat_3248[2]}} | array_update_3251[20] & {32{concat_3248[3]}} | array_update_3252[20] & {32{concat_3248[4]}};
  assign regs__2[21] = array_update_3249[21] & {32{concat_3248[0]}} | regs_unflattened[21] & {32{concat_3248[1]}} | array_update_3250[21] & {32{concat_3248[2]}} | array_update_3251[21] & {32{concat_3248[3]}} | array_update_3252[21] & {32{concat_3248[4]}};
  assign regs__2[22] = array_update_3249[22] & {32{concat_3248[0]}} | regs_unflattened[22] & {32{concat_3248[1]}} | array_update_3250[22] & {32{concat_3248[2]}} | array_update_3251[22] & {32{concat_3248[3]}} | array_update_3252[22] & {32{concat_3248[4]}};
  assign regs__2[23] = array_update_3249[23] & {32{concat_3248[0]}} | regs_unflattened[23] & {32{concat_3248[1]}} | array_update_3250[23] & {32{concat_3248[2]}} | array_update_3251[23] & {32{concat_3248[3]}} | array_update_3252[23] & {32{concat_3248[4]}};
  assign regs__2[24] = array_update_3249[24] & {32{concat_3248[0]}} | regs_unflattened[24] & {32{concat_3248[1]}} | array_update_3250[24] & {32{concat_3248[2]}} | array_update_3251[24] & {32{concat_3248[3]}} | array_update_3252[24] & {32{concat_3248[4]}};
  assign regs__2[25] = array_update_3249[25] & {32{concat_3248[0]}} | regs_unflattened[25] & {32{concat_3248[1]}} | array_update_3250[25] & {32{concat_3248[2]}} | array_update_3251[25] & {32{concat_3248[3]}} | array_update_3252[25] & {32{concat_3248[4]}};
  assign regs__2[26] = array_update_3249[26] & {32{concat_3248[0]}} | regs_unflattened[26] & {32{concat_3248[1]}} | array_update_3250[26] & {32{concat_3248[2]}} | array_update_3251[26] & {32{concat_3248[3]}} | array_update_3252[26] & {32{concat_3248[4]}};
  assign regs__2[27] = array_update_3249[27] & {32{concat_3248[0]}} | regs_unflattened[27] & {32{concat_3248[1]}} | array_update_3250[27] & {32{concat_3248[2]}} | array_update_3251[27] & {32{concat_3248[3]}} | array_update_3252[27] & {32{concat_3248[4]}};
  assign regs__2[28] = array_update_3249[28] & {32{concat_3248[0]}} | regs_unflattened[28] & {32{concat_3248[1]}} | array_update_3250[28] & {32{concat_3248[2]}} | array_update_3251[28] & {32{concat_3248[3]}} | array_update_3252[28] & {32{concat_3248[4]}};
  assign regs__2[29] = array_update_3249[29] & {32{concat_3248[0]}} | regs_unflattened[29] & {32{concat_3248[1]}} | array_update_3250[29] & {32{concat_3248[2]}} | array_update_3251[29] & {32{concat_3248[3]}} | array_update_3252[29] & {32{concat_3248[4]}};
  assign regs__2[30] = array_update_3249[30] & {32{concat_3248[0]}} | regs_unflattened[30] & {32{concat_3248[1]}} | array_update_3250[30] & {32{concat_3248[2]}} | array_update_3251[30] & {32{concat_3248[3]}} | array_update_3252[30] & {32{concat_3248[4]}};
  assign regs__2[31] = array_update_3249[31] & {32{concat_3248[0]}} | regs_unflattened[31] & {32{concat_3248[1]}} | array_update_3250[31] & {32{concat_3248[2]}} | array_update_3251[31] & {32{concat_3248[3]}} | array_update_3252[31] & {32{concat_3248[4]}};
  assign concat_3268 = {and_3193[2:0], opcode__3 != S_CLASS__1 | and_3193[3]};
  assign array_update_3269[0] = add_3257 == 32'h0000_0000 ? array_index_3005[7:0] : dmem__5[0];
  assign array_update_3269[1] = add_3257 == 32'h0000_0001 ? array_index_3005[7:0] : dmem__5[1];
  assign array_update_3269[2] = add_3257 == 32'h0000_0002 ? array_index_3005[7:0] : dmem__5[2];
  assign array_update_3269[3] = add_3257 == 32'h0000_0003 ? array_index_3005[7:0] : dmem__5[3];
  assign array_update_3269[4] = add_3257 == 32'h0000_0004 ? array_index_3005[7:0] : dmem__5[4];
  assign array_update_3269[5] = add_3257 == 32'h0000_0005 ? array_index_3005[7:0] : dmem__5[5];
  assign array_update_3269[6] = add_3257 == 32'h0000_0006 ? array_index_3005[7:0] : dmem__5[6];
  assign array_update_3269[7] = add_3257 == 32'h0000_0007 ? array_index_3005[7:0] : dmem__5[7];
  assign array_update_3269[8] = add_3257 == 32'h0000_0008 ? array_index_3005[7:0] : dmem__5[8];
  assign array_update_3269[9] = add_3257 == 32'h0000_0009 ? array_index_3005[7:0] : dmem__5[9];
  assign array_update_3269[10] = add_3257 == 32'h0000_000a ? array_index_3005[7:0] : dmem__5[10];
  assign array_update_3269[11] = add_3257 == 32'h0000_000b ? array_index_3005[7:0] : dmem__5[11];
  assign array_update_3269[12] = add_3257 == 32'h0000_000c ? array_index_3005[7:0] : dmem__5[12];
  assign array_update_3269[13] = add_3257 == 32'h0000_000d ? array_index_3005[7:0] : dmem__5[13];
  assign array_update_3269[14] = add_3257 == 32'h0000_000e ? array_index_3005[7:0] : dmem__5[14];
  assign array_update_3269[15] = add_3257 == 32'h0000_000f ? array_index_3005[7:0] : dmem__5[15];
  assign array_update_3270[0] = add_3196 == 32'h0000_0000 ? array_index_3005[7:0] : dmem__6[0];
  assign array_update_3270[1] = add_3196 == 32'h0000_0001 ? array_index_3005[7:0] : dmem__6[1];
  assign array_update_3270[2] = add_3196 == 32'h0000_0002 ? array_index_3005[7:0] : dmem__6[2];
  assign array_update_3270[3] = add_3196 == 32'h0000_0003 ? array_index_3005[7:0] : dmem__6[3];
  assign array_update_3270[4] = add_3196 == 32'h0000_0004 ? array_index_3005[7:0] : dmem__6[4];
  assign array_update_3270[5] = add_3196 == 32'h0000_0005 ? array_index_3005[7:0] : dmem__6[5];
  assign array_update_3270[6] = add_3196 == 32'h0000_0006 ? array_index_3005[7:0] : dmem__6[6];
  assign array_update_3270[7] = add_3196 == 32'h0000_0007 ? array_index_3005[7:0] : dmem__6[7];
  assign array_update_3270[8] = add_3196 == 32'h0000_0008 ? array_index_3005[7:0] : dmem__6[8];
  assign array_update_3270[9] = add_3196 == 32'h0000_0009 ? array_index_3005[7:0] : dmem__6[9];
  assign array_update_3270[10] = add_3196 == 32'h0000_000a ? array_index_3005[7:0] : dmem__6[10];
  assign array_update_3270[11] = add_3196 == 32'h0000_000b ? array_index_3005[7:0] : dmem__6[11];
  assign array_update_3270[12] = add_3196 == 32'h0000_000c ? array_index_3005[7:0] : dmem__6[12];
  assign array_update_3270[13] = add_3196 == 32'h0000_000d ? array_index_3005[7:0] : dmem__6[13];
  assign array_update_3270[14] = add_3196 == 32'h0000_000e ? array_index_3005[7:0] : dmem__6[14];
  assign array_update_3270[15] = add_3196 == 32'h0000_000f ? array_index_3005[7:0] : dmem__6[15];
  assign array_update_3271[0] = add_3161 == 32'h0000_0000 ? array_index_3005[7:0] : dmem_unflattened[0];
  assign array_update_3271[1] = add_3161 == 32'h0000_0001 ? array_index_3005[7:0] : dmem_unflattened[1];
  assign array_update_3271[2] = add_3161 == 32'h0000_0002 ? array_index_3005[7:0] : dmem_unflattened[2];
  assign array_update_3271[3] = add_3161 == 32'h0000_0003 ? array_index_3005[7:0] : dmem_unflattened[3];
  assign array_update_3271[4] = add_3161 == 32'h0000_0004 ? array_index_3005[7:0] : dmem_unflattened[4];
  assign array_update_3271[5] = add_3161 == 32'h0000_0005 ? array_index_3005[7:0] : dmem_unflattened[5];
  assign array_update_3271[6] = add_3161 == 32'h0000_0006 ? array_index_3005[7:0] : dmem_unflattened[6];
  assign array_update_3271[7] = add_3161 == 32'h0000_0007 ? array_index_3005[7:0] : dmem_unflattened[7];
  assign array_update_3271[8] = add_3161 == 32'h0000_0008 ? array_index_3005[7:0] : dmem_unflattened[8];
  assign array_update_3271[9] = add_3161 == 32'h0000_0009 ? array_index_3005[7:0] : dmem_unflattened[9];
  assign array_update_3271[10] = add_3161 == 32'h0000_000a ? array_index_3005[7:0] : dmem_unflattened[10];
  assign array_update_3271[11] = add_3161 == 32'h0000_000b ? array_index_3005[7:0] : dmem_unflattened[11];
  assign array_update_3271[12] = add_3161 == 32'h0000_000c ? array_index_3005[7:0] : dmem_unflattened[12];
  assign array_update_3271[13] = add_3161 == 32'h0000_000d ? array_index_3005[7:0] : dmem_unflattened[13];
  assign array_update_3271[14] = add_3161 == 32'h0000_000e ? array_index_3005[7:0] : dmem_unflattened[14];
  assign array_update_3271[15] = add_3161 == 32'h0000_000f ? array_index_3005[7:0] : dmem_unflattened[15];
  assign pc__3 = {add_3073 & {30{concat_3222[0]}} | add_3200[31:2] & {30{concat_3222[1]}} | pc[31:2] & {30{concat_3222[2]}} | sel_3201[31:2] & {30{concat_3222[3]}} | sel_3202[31:2] & {30{concat_3222[4]}} | sel_3203[31:2] & {30{concat_3222[5]}} | sel_3204[31:2] & {30{concat_3222[6]}} | sel_3205[31:2] & {30{concat_3222[7]}} | sel_3206[31:2] & {30{concat_3222[8]}} | add_3207[30:1] & {30{concat_3222[9]}}, pc[1] & concat_3231[0] | add_3200[1] & concat_3231[1] | sel_3201[1] & concat_3231[2] | sel_3202[1] & concat_3231[3] | sel_3203[1] & concat_3231[4] | sel_3204[1] & concat_3231[5] | sel_3205[1] & concat_3231[6] | sel_3206[1] & concat_3231[7] | add_3207[0] & concat_3231[8], pc[0] & concat_3241[0] | sel_3201[0] & concat_3241[1] | sel_3202[0] & concat_3241[2] | sel_3203[0] & concat_3241[3] | sel_3204[0] & concat_3241[4] | sel_3205[0] & concat_3241[5] | sel_3206[0] & concat_3241[6]};
  assign array_update_3277[0] = 32'h0000_0000;
  assign array_update_3277[1] = regs__2[1];
  assign array_update_3277[2] = regs__2[2];
  assign array_update_3277[3] = regs__2[3];
  assign array_update_3277[4] = regs__2[4];
  assign array_update_3277[5] = regs__2[5];
  assign array_update_3277[6] = regs__2[6];
  assign array_update_3277[7] = regs__2[7];
  assign array_update_3277[8] = regs__2[8];
  assign array_update_3277[9] = regs__2[9];
  assign array_update_3277[10] = regs__2[10];
  assign array_update_3277[11] = regs__2[11];
  assign array_update_3277[12] = regs__2[12];
  assign array_update_3277[13] = regs__2[13];
  assign array_update_3277[14] = regs__2[14];
  assign array_update_3277[15] = regs__2[15];
  assign array_update_3277[16] = regs__2[16];
  assign array_update_3277[17] = regs__2[17];
  assign array_update_3277[18] = regs__2[18];
  assign array_update_3277[19] = regs__2[19];
  assign array_update_3277[20] = regs__2[20];
  assign array_update_3277[21] = regs__2[21];
  assign array_update_3277[22] = regs__2[22];
  assign array_update_3277[23] = regs__2[23];
  assign array_update_3277[24] = regs__2[24];
  assign array_update_3277[25] = regs__2[25];
  assign array_update_3277[26] = regs__2[26];
  assign array_update_3277[27] = regs__2[27];
  assign array_update_3277[28] = regs__2[28];
  assign array_update_3277[29] = regs__2[29];
  assign array_update_3277[30] = regs__2[30];
  assign array_update_3277[31] = regs__2[31];
  assign dmem__2[0] = dmem_unflattened[0] & {8{concat_3268[0]}} | array_update_3269[0] & {8{concat_3268[1]}} | array_update_3270[0] & {8{concat_3268[2]}} | array_update_3271[0] & {8{concat_3268[3]}};
  assign dmem__2[1] = dmem_unflattened[1] & {8{concat_3268[0]}} | array_update_3269[1] & {8{concat_3268[1]}} | array_update_3270[1] & {8{concat_3268[2]}} | array_update_3271[1] & {8{concat_3268[3]}};
  assign dmem__2[2] = dmem_unflattened[2] & {8{concat_3268[0]}} | array_update_3269[2] & {8{concat_3268[1]}} | array_update_3270[2] & {8{concat_3268[2]}} | array_update_3271[2] & {8{concat_3268[3]}};
  assign dmem__2[3] = dmem_unflattened[3] & {8{concat_3268[0]}} | array_update_3269[3] & {8{concat_3268[1]}} | array_update_3270[3] & {8{concat_3268[2]}} | array_update_3271[3] & {8{concat_3268[3]}};
  assign dmem__2[4] = dmem_unflattened[4] & {8{concat_3268[0]}} | array_update_3269[4] & {8{concat_3268[1]}} | array_update_3270[4] & {8{concat_3268[2]}} | array_update_3271[4] & {8{concat_3268[3]}};
  assign dmem__2[5] = dmem_unflattened[5] & {8{concat_3268[0]}} | array_update_3269[5] & {8{concat_3268[1]}} | array_update_3270[5] & {8{concat_3268[2]}} | array_update_3271[5] & {8{concat_3268[3]}};
  assign dmem__2[6] = dmem_unflattened[6] & {8{concat_3268[0]}} | array_update_3269[6] & {8{concat_3268[1]}} | array_update_3270[6] & {8{concat_3268[2]}} | array_update_3271[6] & {8{concat_3268[3]}};
  assign dmem__2[7] = dmem_unflattened[7] & {8{concat_3268[0]}} | array_update_3269[7] & {8{concat_3268[1]}} | array_update_3270[7] & {8{concat_3268[2]}} | array_update_3271[7] & {8{concat_3268[3]}};
  assign dmem__2[8] = dmem_unflattened[8] & {8{concat_3268[0]}} | array_update_3269[8] & {8{concat_3268[1]}} | array_update_3270[8] & {8{concat_3268[2]}} | array_update_3271[8] & {8{concat_3268[3]}};
  assign dmem__2[9] = dmem_unflattened[9] & {8{concat_3268[0]}} | array_update_3269[9] & {8{concat_3268[1]}} | array_update_3270[9] & {8{concat_3268[2]}} | array_update_3271[9] & {8{concat_3268[3]}};
  assign dmem__2[10] = dmem_unflattened[10] & {8{concat_3268[0]}} | array_update_3269[10] & {8{concat_3268[1]}} | array_update_3270[10] & {8{concat_3268[2]}} | array_update_3271[10] & {8{concat_3268[3]}};
  assign dmem__2[11] = dmem_unflattened[11] & {8{concat_3268[0]}} | array_update_3269[11] & {8{concat_3268[1]}} | array_update_3270[11] & {8{concat_3268[2]}} | array_update_3271[11] & {8{concat_3268[3]}};
  assign dmem__2[12] = dmem_unflattened[12] & {8{concat_3268[0]}} | array_update_3269[12] & {8{concat_3268[1]}} | array_update_3270[12] & {8{concat_3268[2]}} | array_update_3271[12] & {8{concat_3268[3]}};
  assign dmem__2[13] = dmem_unflattened[13] & {8{concat_3268[0]}} | array_update_3269[13] & {8{concat_3268[1]}} | array_update_3270[13] & {8{concat_3268[2]}} | array_update_3271[13] & {8{concat_3268[3]}};
  assign dmem__2[14] = dmem_unflattened[14] & {8{concat_3268[0]}} | array_update_3269[14] & {8{concat_3268[1]}} | array_update_3270[14] & {8{concat_3268[2]}} | array_update_3271[14] & {8{concat_3268[3]}};
  assign dmem__2[15] = dmem_unflattened[15] & {8{concat_3268[0]}} | array_update_3269[15] & {8{concat_3268[1]}} | array_update_3270[15] & {8{concat_3268[2]}} | array_update_3271[15] & {8{concat_3268[3]}};
  assign out = {pc__3, {array_update_3277[31], array_update_3277[30], array_update_3277[29], array_update_3277[28], array_update_3277[27], array_update_3277[26], array_update_3277[25], array_update_3277[24], array_update_3277[23], array_update_3277[22], array_update_3277[21], array_update_3277[20], array_update_3277[19], array_update_3277[18], array_update_3277[17], array_update_3277[16], array_update_3277[15], array_update_3277[14], array_update_3277[13], array_update_3277[12], array_update_3277[11], array_update_3277[10], array_update_3277[9], array_update_3277[8], array_update_3277[7], array_update_3277[6], array_update_3277[5], array_update_3277[4], array_update_3277[3], array_update_3277[2], array_update_3277[1], array_update_3277[0]}, {dmem__2[15], dmem__2[14], dmem__2[13], dmem__2[12], dmem__2[11], dmem__2[10], dmem__2[9], dmem__2[8], dmem__2[7], dmem__2[6], dmem__2[5], dmem__2[4], dmem__2[3], dmem__2[2], dmem__2[1], dmem__2[0]}};
endmodule
